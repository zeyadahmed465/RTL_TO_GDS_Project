module DLY2X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX3M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI32X2M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22X8M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X3M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX14M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY1X4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module MX2X8M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX1M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFSX2M (
	SN, 
	SI, 
	SE, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX12M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX4M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX2M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2XLM (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI22XLM (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI222XLM (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA22X2M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32XLM (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XNOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFXLM (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX1M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX4M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX8M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X3M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X12M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2XLM (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI33X2M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Sat Sep 23 17:42:53 2023
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN6_RST;
   wire FE_PHN5_RST;
   wire FE_PHN3_scan_reset;
   wire FE_PHN0_scan_reset;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC6_RST (
	.Y(FE_PHN6_RST),
	.A(FE_PHN5_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC5_RST (
	.Y(FE_PHN5_RST),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_scan_reset (
	.Y(FE_PHN3_scan_reset),
	.A(FE_PHN0_scan_reset), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_scan_reset (
	.Y(FE_PHN0_scan_reset),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN3_scan_reset),
	.A(FE_PHN6_RST), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_0 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \sync_reg[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \sync_reg_reg[1]  (
	.SI(\sync_reg[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\sync_reg[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN4_scan_reset;
   wire FE_PHN2_scan_reset;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC4_scan_reset (
	.Y(FE_PHN4_scan_reset),
	.A(FE_PHN2_scan_reset), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_reset (
	.Y(FE_PHN2_scan_reset),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN4_scan_reset),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_1 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \sync_reg[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \sync_reg_reg[1]  (
	.SI(\sync_reg[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\sync_reg[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN1_scan_reset;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC1_scan_reset (
	.Y(FE_PHN1_scan_reset),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN1_scan_reset),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_test_1 (
	CLK, 
	RST, 
	unsync_bus, 
	bus_enable, 
	sync_bus, 
	enable_pulse_d, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] unsync_bus;
   input bus_enable;
   output [7:0] sync_bus;
   output enable_pulse_d;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire enable_flop;
   wire n1;
   wire n4;
   wire n6;
   wire n8;
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n23;
   wire [1:0] sync_reg;

   assign test_so = sync_reg[1] ;

   // Module instantiations
   SDFFRQX2M enable_flop_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(enable_flop),
	.D(sync_reg[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[7]),
	.D(n18),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[5]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[6]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[4]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[3]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[1]),
	.D(n6),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_d_reg (
	.SI(enable_flop),
	.SE(test_se),
	.RN(RST),
	.Q(enable_pulse_d),
	.D(n23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(sync_bus[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[2]),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(enable_pulse_d),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[0]),
	.D(n4),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0]  (
	.SI(sync_bus[7]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_reg[0]),
	.D(bus_enable),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \sync_reg_reg[1]  (
	.SI(sync_reg[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_reg[1]),
	.D(sync_reg[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n23),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U5 (
	.Y(n1),
	.B(sync_reg[1]),
	.AN(enable_flop), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n4),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(n23),
	.A0(unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n6),
	.B1(n1),
	.B0(sync_bus[1]),
	.A1(n23),
	.A0(unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n8),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(n23),
	.A0(unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n10),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(n23),
	.A0(unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n12),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(n23),
	.A0(unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n14),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(n23),
	.A0(unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n16),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(n23),
	.A0(unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n18),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(n23),
	.A0(unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_0 (
	i_ref_clk, 
	i_rst, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	UART_CLK_M__L6_N1, 
	UART_CLK_M__L7_N1, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input UART_CLK_M__L6_N1;
   input UART_CLK_M__L7_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN8_div_clk__Exclude_0_NET;
   wire div_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire N2;
   wire div_clk;
   wire odd_edge_tog;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n3;
   wire n4;
   wire n5;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire [6:0] count;
   wire [6:0] edge_flip_half;

   assign test_so = odd_edge_tog ;

   // Module instantiations
   DLY2X1M FE_PHC8_div_clk__Exclude_0_NET (
	.Y(FE_PHN8_div_clk__Exclude_0_NET),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M div_clk__Exclude_0 (
	.Y(div_clk__Exclude_0_NET),
	.A(div_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[6]  (
	.SI(count[5]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[6]),
	.D(n28),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[0]),
	.D(n34),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[5]  (
	.SI(count[4]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[5]),
	.D(n29),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[4]  (
	.SI(count[3]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[4]),
	.D(n30),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[3]  (
	.SI(count[2]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[3]),
	.D(n31),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(count[1]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[2]),
	.D(n32),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[1]),
	.D(n33),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M odd_edge_tog_reg (
	.SN(i_rst),
	.SI(FE_PHN8_div_clk__Exclude_0_NET),
	.SE(test_se),
	.Q(odd_edge_tog),
	.D(n26),
	.CK(UART_CLK_M__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M div_clk_reg (
	.SI(count[6]),
	.SE(test_se),
	.RN(i_rst),
	.Q(div_clk),
	.D(n27),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U11 (
	.Y(n3),
	.B(i_div_ratio[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U15 (
	.Y(n18),
	.B(HTIE_LTIEHI_NET),
	.AN(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n17),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U17 (
	.Y(o_div_clk),
	.S0(N2),
	.B(div_clk),
	.A(UART_CLK_M__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U18 (
	.Y(edge_flip_half[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U19 (
	.Y(edge_flip_half[1]),
	.B0(n3),
	.A1N(i_div_ratio[2]),
	.A0N(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U20 (
	.Y(n4),
	.B(i_div_ratio[3]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U21 (
	.Y(edge_flip_half[2]),
	.B0(n4),
	.A1N(i_div_ratio[3]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U22 (
	.Y(n5),
	.B(i_div_ratio[4]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U23 (
	.Y(edge_flip_half[3]),
	.B0(n5),
	.A1(i_div_ratio[4]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U24 (
	.Y(n15),
	.B(n17),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U25 (
	.Y(edge_flip_half[4]),
	.B0(n15),
	.A1(n17),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U26 (
	.Y(edge_flip_half[5]),
	.B(n15),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U27 (
	.Y(n16),
	.B(n15),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U28 (
	.Y(edge_flip_half[6]),
	.B(n16),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U29 (
	.Y(n34),
	.B1(n19),
	.B0(N16),
	.A1(count[0]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U30 (
	.Y(n33),
	.B1(n19),
	.B0(N17),
	.A1(count[1]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U31 (
	.Y(n32),
	.B1(n19),
	.B0(N18),
	.A1(count[2]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n31),
	.B1(n19),
	.B0(N19),
	.A1(count[3]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U33 (
	.Y(n30),
	.B1(n19),
	.B0(N20),
	.A1(count[4]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U34 (
	.Y(n29),
	.B1(n19),
	.B0(N21),
	.A1(count[5]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U35 (
	.Y(n28),
	.B1(n19),
	.B0(N22),
	.A1(count[6]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U36 (
	.Y(n19),
	.C(N2),
	.B(n21),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n27),
	.B(n22),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U38 (
	.Y(n22),
	.B0(n18),
	.A1(n20),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U39 (
	.Y(n20),
	.B(i_div_ratio[0]),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U40 (
	.Y(n26),
	.B(n24),
	.A(odd_edge_tog), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U41 (
	.Y(n24),
	.B(n18),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U42 (
	.Y(n21),
	.B(i_div_ratio[0]),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U43 (
	.Y(n25),
	.S0(odd_edge_tog),
	.B(n23),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U44 (
	.Y(n23),
	.D(n39),
	.C(n38),
	.B(n37),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n39),
	.D(n43),
	.C(n42),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n43),
	.B(count[2]),
	.A(edge_flip_half[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n42),
	.B(count[1]),
	.A(edge_flip_half[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n41),
	.B(count[0]),
	.A(edge_flip_half[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n40),
	.B(count[6]),
	.A(edge_flip_half[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n38),
	.B(edge_flip_half[4]),
	.A(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U51 (
	.Y(n37),
	.B(edge_flip_half[5]),
	.A(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U52 (
	.Y(n36),
	.B(edge_flip_half[3]),
	.A(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U53 (
	.Y(n35),
	.D(n47),
	.C(n46),
	.B(n45),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U54 (
	.Y(n47),
	.D(n51),
	.C(n50),
	.B(n49),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n51),
	.B(count[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n50),
	.B(count[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n49),
	.B(count[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n48),
	.B(count[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U59 (
	.Y(n46),
	.B(i_div_ratio[5]),
	.A(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U60 (
	.Y(n45),
	.B(i_div_ratio[6]),
	.A(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U61 (
	.Y(n44),
	.B(i_div_ratio[4]),
	.A(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U62 (
	.Y(N2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U63 (
	.Y(n52),
	.D(i_div_ratio[1]),
	.C(i_div_ratio[3]),
	.B(i_div_ratio[2]),
	.AN(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U64 (
	.Y(n53),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_0_DW01_inc_0 add_49 (
	.A({ count[6],
		count[5],
		count[4],
		count[3],
		count[2],
		count[1],
		count[0] }),
	.SUM({ N22,
		N21,
		N20,
		N19,
		N18,
		N17,
		N16 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_1 (
	i_ref_clk, 
	i_rst, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	UART_CLK_M__L6_N2, 
	UART_CLK_M__L7_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input UART_CLK_M__L6_N2;
   input UART_CLK_M__L7_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_div_clk__Exclude_0_NET;
   wire div_clk__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N2;
   wire div_clk;
   wire odd_edge_tog;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire n3;
   wire n4;
   wire n5;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n74;
   wire n75;
   wire [6:0] count;
   wire [6:0] edge_flip_half;

   assign test_so = odd_edge_tog ;

   // Module instantiations
   DLY2X1M FE_PHC7_div_clk__Exclude_0_NET (
	.Y(FE_PHN7_div_clk__Exclude_0_NET),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M div_clk__Exclude_0 (
	.Y(div_clk__Exclude_0_NET),
	.A(div_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[5]  (
	.SI(count[4]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[5]),
	.D(n59),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[4]  (
	.SI(count[3]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[4]),
	.D(n58),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[3]  (
	.SI(count[2]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[3]),
	.D(n57),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[6]  (
	.SI(count[5]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[6]),
	.D(n60),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[0]),
	.D(n54),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(count[1]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[2]),
	.D(n56),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(test_se),
	.RN(i_rst),
	.Q(count[1]),
	.D(n55),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M div_clk_reg (
	.SI(count[6]),
	.SE(test_se),
	.RN(i_rst),
	.Q(div_clk),
	.D(n61),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U11 (
	.Y(n18),
	.B(HTIE_LTIEHI_NET),
	.AN(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n17),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U16 (
	.Y(n3),
	.B(LTIE_LTIELO_NET),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U17 (
	.Y(o_div_clk),
	.S0(N2),
	.B(div_clk),
	.A(UART_CLK_M__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U18 (
	.Y(edge_flip_half[0]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U19 (
	.Y(edge_flip_half[1]),
	.B0(n3),
	.A1N(HTIE_LTIEHI_NET),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U20 (
	.Y(n4),
	.B(LTIE_LTIELO_NET),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U21 (
	.Y(edge_flip_half[2]),
	.B0(n4),
	.A1N(LTIE_LTIELO_NET),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U22 (
	.Y(n5),
	.B(LTIE_LTIELO_NET),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U23 (
	.Y(edge_flip_half[3]),
	.B0(n5),
	.A1(LTIE_LTIELO_NET),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U24 (
	.Y(n15),
	.B(n17),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U25 (
	.Y(edge_flip_half[4]),
	.B0(n15),
	.A1(n17),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U26 (
	.Y(edge_flip_half[5]),
	.B(n15),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U27 (
	.Y(n16),
	.B(n15),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U28 (
	.Y(edge_flip_half[6]),
	.B(n16),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U29 (
	.Y(n54),
	.B1(n19),
	.B0(N16),
	.A1(count[0]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U30 (
	.Y(n55),
	.B1(n19),
	.B0(N17),
	.A1(count[1]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U31 (
	.Y(n56),
	.B1(n19),
	.B0(N18),
	.A1(count[2]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n57),
	.B1(n19),
	.B0(N19),
	.A1(count[3]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U33 (
	.Y(n58),
	.B1(n19),
	.B0(N20),
	.A1(count[4]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U34 (
	.Y(n59),
	.B1(n19),
	.B0(N21),
	.A1(count[5]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U35 (
	.Y(n60),
	.B1(n19),
	.B0(N22),
	.A1(count[6]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U36 (
	.Y(n19),
	.C(N2),
	.B(n21),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n61),
	.B(n22),
	.A(div_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U38 (
	.Y(n22),
	.B0(n18),
	.A1(n20),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U39 (
	.Y(n20),
	.B(LTIE_LTIELO_NET),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U40 (
	.Y(n62),
	.B(n24),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U41 (
	.Y(n24),
	.B(n18),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U42 (
	.Y(n21),
	.B(LTIE_LTIELO_NET),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U43 (
	.Y(n25),
	.S0(n75),
	.B(n23),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U44 (
	.Y(n23),
	.D(n39),
	.C(n38),
	.B(n37),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n39),
	.D(n43),
	.C(n42),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U46 (
	.Y(n43),
	.B(count[2]),
	.A(edge_flip_half[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n42),
	.B(count[1]),
	.A(edge_flip_half[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n41),
	.B(count[0]),
	.A(edge_flip_half[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n40),
	.B(count[6]),
	.A(edge_flip_half[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n38),
	.B(edge_flip_half[4]),
	.A(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U51 (
	.Y(n37),
	.B(edge_flip_half[5]),
	.A(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U52 (
	.Y(n36),
	.B(edge_flip_half[3]),
	.A(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U53 (
	.Y(n35),
	.D(n47),
	.C(n46),
	.B(n45),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U54 (
	.Y(n47),
	.D(n51),
	.C(n50),
	.B(n49),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n51),
	.B(count[2]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n50),
	.B(count[1]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n49),
	.B(count[0]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n48),
	.B(count[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U59 (
	.Y(n46),
	.B(LTIE_LTIELO_NET),
	.A(count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U60 (
	.Y(n45),
	.B(LTIE_LTIELO_NET),
	.A(count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U61 (
	.Y(n44),
	.B(LTIE_LTIELO_NET),
	.A(count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U62 (
	.Y(N2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U63 (
	.Y(n52),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(HTIE_LTIEHI_NET),
	.AN(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U64 (
	.Y(n53),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U66 (
	.Y(n75),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_1_DW01_inc_0 add_49 (
	.A({ count[6],
		count[5],
		count[4],
		count[3],
		count[2],
		count[1],
		count[0] }),
	.SUM({ N22,
		N21,
		N20,
		N19,
		N18,
		N17,
		N16 }), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSX2M odd_edge_tog_reg (
	.SN(i_rst),
	.SI(FE_PHN7_div_clk__Exclude_0_NET),
	.SE(test_se),
	.QN(n74),
	.Q(odd_edge_tog),
	.D(n62),
	.CK(UART_CLK_M__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_GATE (
	CLK_EN, 
	CLK, 
	GATED_CLK, 
	VDD, 
	VSS);
   input CLK_EN;
   input CLK;
   output GATED_CLK;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX12M U0_TLATNCAX12M (
	.ECK(GATED_CLK),
	.E(CLK_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module REG_FILE_test_1 (
	WrData, 
	Address, 
	WrEn, 
	RdEn, 
	CLK, 
	RST, 
	RdData, 
	RdData_VLD, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] WrData;
   input [3:0] Address;
   input WrEn;
   input RdEn;
   input CLK;
   input RST;
   output [7:0] RdData;
   output RdData_VLD;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN10_Op_B_7_;
   wire FE_OFN9_Op_B_1_;
   wire FE_OFN8_Op_A_6_;
   wire FE_OFN7_Op_A_5_;
   wire FE_OFN6_Op_B_6_;
   wire FE_OFN5_Op_A_7_;
   wire FE_OFN2_SYNC_REF_RST_M;
   wire FE_OFN1_SYNC_REF_RST_M;
   wire \Reg_File[13][7] ;
   wire \Reg_File[13][6] ;
   wire \Reg_File[13][5] ;
   wire \Reg_File[13][4] ;
   wire \Reg_File[13][3] ;
   wire \Reg_File[13][2] ;
   wire \Reg_File[13][1] ;
   wire \Reg_File[13][0] ;
   wire \Reg_File[12][7] ;
   wire \Reg_File[12][6] ;
   wire \Reg_File[12][5] ;
   wire \Reg_File[12][4] ;
   wire \Reg_File[12][3] ;
   wire \Reg_File[12][2] ;
   wire \Reg_File[12][1] ;
   wire \Reg_File[12][0] ;
   wire \Reg_File[9][7] ;
   wire \Reg_File[9][6] ;
   wire \Reg_File[9][5] ;
   wire \Reg_File[9][4] ;
   wire \Reg_File[9][3] ;
   wire \Reg_File[9][2] ;
   wire \Reg_File[9][1] ;
   wire \Reg_File[9][0] ;
   wire \Reg_File[8][7] ;
   wire \Reg_File[8][6] ;
   wire \Reg_File[8][5] ;
   wire \Reg_File[8][4] ;
   wire \Reg_File[8][3] ;
   wire \Reg_File[8][2] ;
   wire \Reg_File[8][1] ;
   wire \Reg_File[8][0] ;
   wire \Reg_File[7][7] ;
   wire \Reg_File[7][6] ;
   wire \Reg_File[7][5] ;
   wire \Reg_File[7][4] ;
   wire \Reg_File[7][3] ;
   wire \Reg_File[7][2] ;
   wire \Reg_File[7][1] ;
   wire \Reg_File[7][0] ;
   wire \Reg_File[6][7] ;
   wire \Reg_File[6][6] ;
   wire \Reg_File[6][5] ;
   wire \Reg_File[6][4] ;
   wire \Reg_File[6][3] ;
   wire \Reg_File[6][2] ;
   wire \Reg_File[6][1] ;
   wire \Reg_File[6][0] ;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n186;
   wire n208;
   wire n280;
   wire n290;
   wire n310;
   wire n473;
   wire n476;
   wire n478;
   wire n480;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n563;
   wire n564;
   wire n565;
   wire n566;

   assign test_so1 = \Reg_File[13][6]  ;

   // Module instantiations
   BUFX14M FE_OFC10_Op_B_7_ (
	.Y(REG1[7]),
	.A(FE_OFN10_Op_B_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC9_Op_B_1_ (
	.Y(REG1[1]),
	.A(FE_OFN9_Op_B_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC8_Op_A_6_ (
	.Y(REG0[6]),
	.A(FE_OFN8_Op_A_6_), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M FE_OFC7_Op_A_5_ (
	.Y(REG0[5]),
	.A(FE_OFN7_Op_A_5_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC6_Op_B_6_ (
	.Y(REG1[6]),
	.A(FE_OFN6_Op_B_6_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC5_Op_A_7_ (
	.Y(REG0[7]),
	.A(FE_OFN5_Op_A_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX6M FE_OFC2_SYNC_REF_RST_M (
	.Y(FE_OFN2_SYNC_REF_RST_M),
	.A(FE_OFN1_SYNC_REF_RST_M), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC1_SYNC_REF_RST_M (
	.Y(FE_OFN1_SYNC_REF_RST_M),
	.A(RST), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \Reg_File_reg[1][7]  (
	.SI(REG1[6]),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(FE_OFN10_Op_B_7_),
	.D(n359),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][2]  (
	.SI(REG2[1]),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[2]),
	.D(n362),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][7]  (
	.SI(\Reg_File[6][6] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][7] ),
	.D(n399),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][6]  (
	.SI(\Reg_File[6][5] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][6] ),
	.D(n398),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][5]  (
	.SI(\Reg_File[6][4] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][5] ),
	.D(n397),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][4]  (
	.SI(\Reg_File[6][3] ),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][4] ),
	.D(n396),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][3]  (
	.SI(\Reg_File[6][2] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][3] ),
	.D(n395),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][2]  (
	.SI(\Reg_File[6][1] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][2] ),
	.D(n394),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][1]  (
	.SI(\Reg_File[6][0] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][1] ),
	.D(n393),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[6][0]  (
	.SI(n539),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[6][0] ),
	.D(n392),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[7]  (
	.SI(RdData[6]),
	.SE(n566),
	.RN(RST),
	.Q(RdData[7]),
	.D(n342),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[6]  (
	.SI(RdData[5]),
	.SE(n565),
	.RN(RST),
	.Q(RdData[6]),
	.D(n341),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[5]  (
	.SI(RdData[4]),
	.SE(n564),
	.RN(RST),
	.Q(RdData[5]),
	.D(n340),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[4]  (
	.SI(RdData[3]),
	.SE(n563),
	.RN(RST),
	.Q(RdData[4]),
	.D(n339),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[3]  (
	.SI(RdData[2]),
	.SE(n566),
	.RN(RST),
	.Q(RdData[3]),
	.D(n338),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[2]  (
	.SI(RdData[1]),
	.SE(n565),
	.RN(RST),
	.Q(RdData[2]),
	.D(n337),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[1]  (
	.SI(RdData[0]),
	.SE(n564),
	.RN(RST),
	.Q(RdData[1]),
	.D(n336),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[0]  (
	.SI(RdData_VLD),
	.SE(n563),
	.RN(RST),
	.Q(RdData[0]),
	.D(n335),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][7]  (
	.SI(\Reg_File[7][6] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][7] ),
	.D(n407),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][6]  (
	.SI(\Reg_File[7][5] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][6] ),
	.D(n406),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][5]  (
	.SI(\Reg_File[7][4] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][5] ),
	.D(n405),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][4]  (
	.SI(\Reg_File[7][3] ),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][4] ),
	.D(n404),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][3]  (
	.SI(\Reg_File[7][2] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][3] ),
	.D(n403),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][2]  (
	.SI(\Reg_File[7][1] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][2] ),
	.D(n402),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][1]  (
	.SI(\Reg_File[7][0] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][1] ),
	.D(n401),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[7][0]  (
	.SI(\Reg_File[6][7] ),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[7][0] ),
	.D(n400),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][7]  (
	.SI(test_si3),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[13][7] ),
	.D(n455),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][6]  (
	.SI(\Reg_File[13][5] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[13][6] ),
	.D(n454),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][5]  (
	.SI(\Reg_File[13][4] ),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[13][5] ),
	.D(n453),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][4]  (
	.SI(\Reg_File[13][3] ),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[13][4] ),
	.D(n452),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][3]  (
	.SI(\Reg_File[13][2] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[13][3] ),
	.D(n451),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][2]  (
	.SI(\Reg_File[13][1] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[13][2] ),
	.D(n450),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][1]  (
	.SI(\Reg_File[13][0] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[13][1] ),
	.D(n449),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[13][0]  (
	.SI(\Reg_File[12][7] ),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[13][0] ),
	.D(n448),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][7]  (
	.SI(\Reg_File[9][6] ),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][7] ),
	.D(n423),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][6]  (
	.SI(\Reg_File[9][5] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][6] ),
	.D(n422),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][5]  (
	.SI(\Reg_File[9][4] ),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][5] ),
	.D(n421),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][4]  (
	.SI(\Reg_File[9][3] ),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][4] ),
	.D(n420),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][3]  (
	.SI(\Reg_File[9][2] ),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][3] ),
	.D(n419),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][2]  (
	.SI(\Reg_File[9][1] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][2] ),
	.D(n418),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][1]  (
	.SI(\Reg_File[9][0] ),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][1] ),
	.D(n417),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[9][0]  (
	.SI(\Reg_File[8][7] ),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[9][0] ),
	.D(n416),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][7]  (
	.SI(\Reg_File[12][6] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][7] ),
	.D(n447),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][6]  (
	.SI(\Reg_File[12][5] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][6] ),
	.D(n446),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][5]  (
	.SI(\Reg_File[12][4] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][5] ),
	.D(n445),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][4]  (
	.SI(\Reg_File[12][3] ),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][4] ),
	.D(n444),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][3]  (
	.SI(\Reg_File[12][2] ),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][3] ),
	.D(n443),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][2]  (
	.SI(\Reg_File[12][1] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][2] ),
	.D(n442),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][1]  (
	.SI(\Reg_File[12][0] ),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][1] ),
	.D(n441),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[12][0]  (
	.SI(n523),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(\Reg_File[12][0] ),
	.D(n440),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][7]  (
	.SI(\Reg_File[8][6] ),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][7] ),
	.D(n415),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][6]  (
	.SI(\Reg_File[8][5] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][6] ),
	.D(n414),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][5]  (
	.SI(\Reg_File[8][4] ),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][5] ),
	.D(n413),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][4]  (
	.SI(\Reg_File[8][3] ),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][4] ),
	.D(n412),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][3]  (
	.SI(\Reg_File[8][2] ),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][3] ),
	.D(n411),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][2]  (
	.SI(\Reg_File[8][1] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][2] ),
	.D(n410),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][1]  (
	.SI(\Reg_File[8][0] ),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][1] ),
	.D(n409),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[8][0]  (
	.SI(\Reg_File[7][7] ),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(\Reg_File[8][0] ),
	.D(n408),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][0]  (
	.SI(REG2[7]),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[0]),
	.D(n368),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][1]  (
	.SI(REG2[0]),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[1]),
	.D(n361),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][4]  (
	.SI(REG3[3]),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[4]),
	.D(n372),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \Reg_File_reg[3][2]  (
	.SI(REG3[1]),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[2]),
	.D(n370),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][3]  (
	.SI(test_si2),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[3]),
	.D(n371),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][7]  (
	.SI(n516),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n146),
	.Q(n515),
	.D(n463),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][6]  (
	.SI(n517),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n147),
	.Q(n516),
	.D(n462),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][5]  (
	.SI(n518),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n148),
	.Q(n517),
	.D(n461),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][4]  (
	.SI(n519),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n149),
	.Q(n518),
	.D(n460),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][3]  (
	.SI(n520),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n150),
	.Q(n519),
	.D(n459),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][2]  (
	.SI(n521),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n151),
	.Q(n520),
	.D(n458),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][1]  (
	.SI(n522),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n152),
	.Q(n521),
	.D(n457),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[14][0]  (
	.SI(\Reg_File[13][7] ),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n153),
	.Q(n522),
	.D(n456),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][7]  (
	.SI(n532),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n162),
	.Q(n531),
	.D(n431),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][6]  (
	.SI(n533),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n163),
	.Q(n532),
	.D(n430),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][5]  (
	.SI(n534),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n164),
	.Q(n533),
	.D(n429),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][4]  (
	.SI(n535),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n165),
	.Q(n534),
	.D(n428),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][3]  (
	.SI(n536),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n166),
	.Q(n535),
	.D(n427),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][2]  (
	.SI(n537),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n167),
	.Q(n536),
	.D(n426),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][1]  (
	.SI(n538),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n168),
	.Q(n537),
	.D(n425),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[10][0]  (
	.SI(\Reg_File[9][7] ),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n169),
	.Q(n538),
	.D(n424),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][7]  (
	.SI(n508),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n138),
	.Q(test_so2),
	.D(n471),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][6]  (
	.SI(n509),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n139),
	.Q(n508),
	.D(n470),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][5]  (
	.SI(n510),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n140),
	.Q(n509),
	.D(n469),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][4]  (
	.SI(n511),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n141),
	.Q(n510),
	.D(n468),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][3]  (
	.SI(n512),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n142),
	.Q(n511),
	.D(n467),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][2]  (
	.SI(n513),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n143),
	.Q(n512),
	.D(n466),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][1]  (
	.SI(n514),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n144),
	.Q(n513),
	.D(n465),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[15][0]  (
	.SI(n515),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n145),
	.Q(n514),
	.D(n464),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][6]  (
	.SI(n525),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n155),
	.Q(n524),
	.D(n438),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][5]  (
	.SI(n526),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n156),
	.Q(n525),
	.D(n437),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][4]  (
	.SI(n527),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n157),
	.Q(n526),
	.D(n436),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][3]  (
	.SI(n528),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n158),
	.Q(n527),
	.D(n435),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][2]  (
	.SI(n529),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n159),
	.Q(n528),
	.D(n434),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][1]  (
	.SI(n530),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n160),
	.Q(n529),
	.D(n433),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][0]  (
	.SI(n531),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n161),
	.Q(n530),
	.D(n432),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][7]  (
	.SI(n540),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n170),
	.Q(n539),
	.D(n391),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][6]  (
	.SI(n541),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n171),
	.Q(n540),
	.D(n390),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][5]  (
	.SI(n542),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n172),
	.Q(n541),
	.D(n389),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][4]  (
	.SI(n543),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n173),
	.Q(n542),
	.D(n388),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][3]  (
	.SI(n544),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n174),
	.Q(n543),
	.D(n387),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][2]  (
	.SI(n545),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n175),
	.Q(n544),
	.D(n386),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][1]  (
	.SI(n546),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n176),
	.Q(n545),
	.D(n385),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[5][0]  (
	.SI(n547),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n177),
	.Q(n546),
	.D(n384),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][7]  (
	.SI(n548),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n178),
	.Q(n547),
	.D(n383),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][6]  (
	.SI(n549),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n179),
	.Q(n548),
	.D(n382),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][5]  (
	.SI(n550),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n180),
	.Q(n549),
	.D(n381),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][4]  (
	.SI(n551),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n181),
	.Q(n550),
	.D(n380),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][3]  (
	.SI(n552),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n182),
	.Q(n551),
	.D(n379),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][2]  (
	.SI(n553),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n183),
	.Q(n552),
	.D(n378),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][1]  (
	.SI(n554),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n184),
	.Q(n553),
	.D(n377),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[4][0]  (
	.SI(REG3[7]),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n185),
	.Q(n554),
	.D(n376),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][1]  (
	.SI(REG3[0]),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[1]),
	.D(n369),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][3]  (
	.SI(REG2[2]),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[3]),
	.D(n363),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \Reg_File_reg[2][0]  (
	.SN(FE_OFN2_SYNC_REF_RST_M),
	.SI(REG1[7]),
	.SE(n563),
	.Q(REG2[0]),
	.D(n360),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][4]  (
	.SI(REG2[3]),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[4]),
	.D(n364),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RdData_VLD_reg (
	.SI(test_si1),
	.SE(n566),
	.RN(RST),
	.Q(RdData_VLD),
	.D(n343),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][7]  (
	.SI(REG2[6]),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[7]),
	.D(n367),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[2][6]  (
	.SI(REG2[5]),
	.SE(n563),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG2[6]),
	.D(n366),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][6]  (
	.SI(REG3[5]),
	.SE(n566),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[6]),
	.D(n374),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Reg_File_reg[3][7]  (
	.SI(REG3[6]),
	.SE(n565),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.Q(REG3[7]),
	.D(n375),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX4M \Reg_File_reg[1][2]  (
	.SI(REG1[1]),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n191),
	.Q(n558),
	.D(n354),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M \Reg_File_reg[3][5]  (
	.SN(FE_OFN1_SYNC_REF_RST_M),
	.SI(REG3[4]),
	.SE(n566),
	.Q(REG3[5]),
	.D(n373),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[11][7]  (
	.SI(n524),
	.SE(n564),
	.RN(FE_OFN1_SYNC_REF_RST_M),
	.QN(n154),
	.Q(n523),
	.D(n439),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \Reg_File_reg[1][1]  (
	.SI(REG1[0]),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(FE_OFN9_Op_B_1_),
	.D(n353),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[0][4]  (
	.SI(n198),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n197),
	.Q(REG0[4]),
	.D(n348),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[0][3]  (
	.SI(n199),
	.SE(n566),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n198),
	.Q(REG0[3]),
	.D(n347),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[0][2]  (
	.SI(n200),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n199),
	.Q(REG0[2]),
	.D(n346),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[0][1]  (
	.SI(n201),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n200),
	.Q(REG0[1]),
	.D(n345),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Reg_File_reg[0][0]  (
	.SI(RdData[7]),
	.SE(n563),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.QN(n201),
	.Q(REG0[0]),
	.D(n344),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \Reg_File_reg[0][6]  (
	.SI(REG0[5]),
	.SE(n564),
	.RN(RST),
	.Q(FE_OFN8_Op_A_6_),
	.D(n350),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \Reg_File_reg[0][5]  (
	.SI(n197),
	.SE(n564),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(FE_OFN7_Op_A_5_),
	.D(n349),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M \Reg_File_reg[2][5]  (
	.SN(FE_OFN1_SYNC_REF_RST_M),
	.SI(REG2[4]),
	.SE(n565),
	.Q(REG2[5]),
	.D(n365),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX4M \Reg_File_reg[1][5]  (
	.SI(n556),
	.SE(n566),
	.RN(RST),
	.QN(n188),
	.Q(n555),
	.D(n357),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX4M \Reg_File_reg[1][4]  (
	.SI(n557),
	.SE(n565),
	.RN(RST),
	.QN(n189),
	.Q(n556),
	.D(n356),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX2M \Reg_File_reg[1][3]  (
	.SI(n558),
	.SE(test_se),
	.RN(RST),
	.QN(n190),
	.Q(n557),
	.D(n355),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \Reg_File_reg[1][6]  (
	.SI(n555),
	.SE(n563),
	.RN(RST),
	.Q(FE_OFN6_Op_B_6_),
	.D(n358),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \Reg_File_reg[1][0]  (
	.SI(REG0[7]),
	.SE(n565),
	.RN(FE_OFN2_SYNC_REF_RST_M),
	.Q(n484),
	.D(n352),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \Reg_File_reg[0][7]  (
	.SI(REG0[6]),
	.SE(n564),
	.RN(RST),
	.Q(FE_OFN5_Op_A_7_),
	.D(n351),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U140 (
	.Y(REG1[4]),
	.A(n189), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U141 (
	.Y(REG1[5]),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U142 (
	.Y(n186),
	.B(n492),
	.A(n280), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U143 (
	.Y(REG1[3]),
	.A(n190), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U155 (
	.Y(n208),
	.A(n484), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U156 (
	.Y(REG1[0]),
	.A(n208), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U157 (
	.Y(n352),
	.S0(n186),
	.B(WrData[0]),
	.A(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U158 (
	.Y(n321),
	.B(n233),
	.AN(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U159 (
	.Y(n491),
	.A(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U160 (
	.Y(n488),
	.A(n328), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U161 (
	.Y(n487),
	.A(n329), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U162 (
	.Y(n486),
	.A(n333), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U163 (
	.Y(n485),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U164 (
	.Y(n490),
	.A(n320), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U165 (
	.Y(n489),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n318),
	.B(n493),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n319),
	.B(n495),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n323),
	.B(n493),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n324),
	.B(n495),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U170 (
	.Y(n325),
	.B(n241),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U171 (
	.Y(n327),
	.B(n242),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U172 (
	.Y(n330),
	.B(n241),
	.A(n331), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U173 (
	.Y(n332),
	.B(n242),
	.A(n331), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U174 (
	.Y(n315),
	.B(n241),
	.AN(n280), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U175 (
	.Y(n328),
	.B(n493),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U176 (
	.Y(n329),
	.B(n495),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U177 (
	.Y(n333),
	.B(n493),
	.A(n331), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U178 (
	.Y(n334),
	.B(n495),
	.A(n331), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U179 (
	.Y(n320),
	.B(n241),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U180 (
	.Y(n322),
	.B(n242),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U181 (
	.Y(n492),
	.A(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U182 (
	.Y(n496),
	.A(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U183 (
	.Y(n280),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U184 (
	.Y(n316),
	.B(n235),
	.AN(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U185 (
	.Y(n493),
	.A(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U186 (
	.Y(n495),
	.A(n239), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U187 (
	.Y(n331),
	.B(n229),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U188 (
	.Y(n326),
	.B(n227),
	.A(n314), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U193 (
	.Y(n238),
	.B(n494),
	.A(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U194 (
	.Y(n239),
	.B(Address[0]),
	.A(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U195 (
	.Y(n314),
	.B(RdEn),
	.AN(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U196 (
	.Y(n242),
	.B(Address[1]),
	.A(n494), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U197 (
	.Y(n241),
	.B(Address[1]),
	.A(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U198 (
	.Y(n494),
	.A(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U199 (
	.Y(n226),
	.B(RdEn),
	.AN(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U200 (
	.Y(n499),
	.A(WrData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U201 (
	.Y(n500),
	.A(WrData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U202 (
	.Y(n501),
	.A(WrData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U203 (
	.Y(n502),
	.A(WrData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U204 (
	.Y(n503),
	.A(WrData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U205 (
	.Y(n504),
	.A(WrData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U206 (
	.Y(n229),
	.B(n497),
	.A(n498), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U207 (
	.Y(n227),
	.B(Address[2]),
	.A(n498), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U208 (
	.Y(n235),
	.B(n498),
	.A(n497), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U209 (
	.Y(n233),
	.B(n498),
	.A(Address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U210 (
	.Y(n497),
	.A(Address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U220 (
	.Y(n349),
	.S0(n491),
	.B(WrData[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U221 (
	.Y(n350),
	.S0(n491),
	.B(WrData[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U222 (
	.Y(n354),
	.S0(n186),
	.B(WrData[2]),
	.A(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U223 (
	.Y(n355),
	.S0(n186),
	.B(WrData[3]),
	.A(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U224 (
	.Y(n356),
	.S0(n186),
	.B(WrData[4]),
	.A(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U225 (
	.Y(n357),
	.S0(n186),
	.B(WrData[5]),
	.A(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U226 (
	.Y(n505),
	.A(WrData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U227 (
	.Y(n506),
	.A(WrData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U228 (
	.Y(n498),
	.A(Address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U232 (
	.Y(n307),
	.B1(n235),
	.B0(n309),
	.A1(n233),
	.A0(n308), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U233 (
	.Y(n308),
	.C0(n311),
	.B1(n495),
	.B0(\Reg_File[7][7] ),
	.A1(n493),
	.A0(\Reg_File[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U234 (
	.Y(n311),
	.B1(n178),
	.B0(n496),
	.A1(n170),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n335),
	.B1(n226),
	.B0(n225),
	.A1N(n226),
	.A0N(RdData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U236 (
	.Y(n225),
	.C0(n231),
	.B1(n230),
	.B0(n229),
	.A1(n228),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U237 (
	.Y(n228),
	.C0(n243),
	.B1(n161),
	.B0(n239),
	.A1(n169),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U238 (
	.Y(n230),
	.C0(n240),
	.B1(n145),
	.B0(n239),
	.A1(n153),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n336),
	.B1(n226),
	.B0(n244),
	.A1N(n226),
	.A0N(RdData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U240 (
	.Y(n244),
	.C0(n247),
	.B1(n246),
	.B0(n229),
	.A1(n245),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U241 (
	.Y(n245),
	.C0(n253),
	.B1(n160),
	.B0(n239),
	.A1(n168),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U242 (
	.Y(n246),
	.C0(n252),
	.B1(n144),
	.B0(n239),
	.A1(n152),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n337),
	.B1(n226),
	.B0(n254),
	.A1N(n226),
	.A0N(RdData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U244 (
	.Y(n254),
	.C0(n257),
	.B1(n256),
	.B0(n229),
	.A1(n255),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U245 (
	.Y(n255),
	.C0(n263),
	.B1(n159),
	.B0(n239),
	.A1(n167),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U246 (
	.Y(n256),
	.C0(n262),
	.B1(n143),
	.B0(n239),
	.A1(n151),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n338),
	.B1(n226),
	.B0(n264),
	.A1N(n226),
	.A0N(RdData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U248 (
	.Y(n264),
	.C0(n267),
	.B1(n266),
	.B0(n229),
	.A1(n265),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U249 (
	.Y(n265),
	.C0(n273),
	.B1(n158),
	.B0(n239),
	.A1(n166),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U250 (
	.Y(n266),
	.C0(n272),
	.B1(n142),
	.B0(n239),
	.A1(n150),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n339),
	.B1(n226),
	.B0(n274),
	.A1N(n226),
	.A0N(RdData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U252 (
	.Y(n274),
	.C0(n277),
	.B1(n276),
	.B0(n229),
	.A1(n275),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U253 (
	.Y(n275),
	.C0(n283),
	.B1(n157),
	.B0(n239),
	.A1(n165),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U254 (
	.Y(n276),
	.C0(n282),
	.B1(n141),
	.B0(n239),
	.A1(n149),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n340),
	.B1(n226),
	.B0(n284),
	.A1N(n226),
	.A0N(RdData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U256 (
	.Y(n284),
	.C0(n287),
	.B1(n286),
	.B0(n229),
	.A1(n285),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U257 (
	.Y(n285),
	.C0(n293),
	.B1(n156),
	.B0(n239),
	.A1(n164),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U258 (
	.Y(n286),
	.C0(n292),
	.B1(n140),
	.B0(n239),
	.A1(n148),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n341),
	.B1(n226),
	.B0(n294),
	.A1N(n226),
	.A0N(RdData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221X1M U260 (
	.Y(n294),
	.C0(n297),
	.B1(n296),
	.B0(n229),
	.A1(n295),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U261 (
	.Y(n295),
	.C0(n303),
	.B1(n155),
	.B0(n239),
	.A1(n163),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U262 (
	.Y(n296),
	.C0(n302),
	.B1(n139),
	.B0(n239),
	.A1(n147),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n342),
	.B1(n226),
	.B0(n304),
	.A1N(n226),
	.A0N(RdData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U264 (
	.Y(n304),
	.C0(n307),
	.B1(n306),
	.B0(n229),
	.A1(n305),
	.A0(n227), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U265 (
	.Y(n305),
	.C0(n313),
	.B1(n154),
	.B0(n239),
	.A1(n162),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U266 (
	.Y(n306),
	.C0(n312),
	.B1(n138),
	.B0(n239),
	.A1(n146),
	.A0(n238), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U267 (
	.Y(n297),
	.B1(n235),
	.B0(n299),
	.A1(n233),
	.A0(n298), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U268 (
	.Y(n298),
	.C0(n301),
	.B1(n495),
	.B0(\Reg_File[7][6] ),
	.A1(n493),
	.A0(\Reg_File[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U269 (
	.Y(n301),
	.B1(n179),
	.B0(n496),
	.A1(n171),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U270 (
	.Y(n247),
	.B1(n235),
	.B0(n249),
	.A1(n233),
	.A0(n248), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U271 (
	.Y(n248),
	.C0(n251),
	.B1(n495),
	.B0(\Reg_File[7][1] ),
	.A1(n493),
	.A0(\Reg_File[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U272 (
	.Y(n249),
	.C0(n482),
	.B1(n242),
	.B0(REG1[1]),
	.A1(REG0[1]),
	.A0(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U273 (
	.Y(n251),
	.B1(n184),
	.B0(n496),
	.A1(n176),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U274 (
	.Y(n257),
	.B1(n235),
	.B0(n259),
	.A1(n233),
	.A0(n258), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U275 (
	.Y(n258),
	.C0(n261),
	.B1(n495),
	.B0(\Reg_File[7][2] ),
	.A1(n493),
	.A0(\Reg_File[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U276 (
	.Y(n259),
	.C0(n480),
	.B1(n242),
	.B0(REG1[2]),
	.A1(REG0[2]),
	.A0(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U277 (
	.Y(n261),
	.B1(n183),
	.B0(n496),
	.A1(n175),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U278 (
	.Y(n267),
	.B1(n235),
	.B0(n269),
	.A1(n233),
	.A0(n268), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U279 (
	.Y(n268),
	.C0(n271),
	.B1(n495),
	.B0(\Reg_File[7][3] ),
	.A1(n493),
	.A0(\Reg_File[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U280 (
	.Y(n269),
	.C0(n478),
	.B1(n242),
	.B0(REG1[3]),
	.A1(REG0[3]),
	.A0(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U281 (
	.Y(n271),
	.B1(n182),
	.B0(n496),
	.A1(n174),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U282 (
	.Y(n277),
	.B1(n235),
	.B0(n279),
	.A1(n233),
	.A0(n278), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U283 (
	.Y(n278),
	.C0(n281),
	.B1(n495),
	.B0(\Reg_File[7][4] ),
	.A1(n493),
	.A0(\Reg_File[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U284 (
	.Y(n279),
	.C0(n476),
	.B1(n242),
	.B0(REG1[4]),
	.A1(REG0[4]),
	.A0(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U285 (
	.Y(n281),
	.B1(n181),
	.B0(n496),
	.A1(n173),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U286 (
	.Y(n287),
	.B1(n235),
	.B0(n289),
	.A1(n233),
	.A0(n288), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U287 (
	.Y(n288),
	.C0(n291),
	.B1(n495),
	.B0(\Reg_File[7][5] ),
	.A1(n493),
	.A0(\Reg_File[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U288 (
	.Y(n289),
	.C0(n473),
	.B1(n242),
	.B0(REG1[5]),
	.A1(n241),
	.A0(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U289 (
	.Y(n291),
	.B1(n180),
	.B0(n496),
	.A1(n172),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U290 (
	.Y(n231),
	.B1(n235),
	.B0(n234),
	.A1(n233),
	.A0(n232), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U291 (
	.Y(n232),
	.C0(n237),
	.B1(n495),
	.B0(\Reg_File[7][0] ),
	.A1(n493),
	.A0(\Reg_File[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U292 (
	.Y(n234),
	.C0(n483),
	.B1(n242),
	.B0(REG1[0]),
	.A1(REG0[0]),
	.A0(n241), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U293 (
	.Y(n237),
	.B1(n185),
	.B0(n496),
	.A1(n177),
	.A0(n492), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U294 (
	.Y(n424),
	.B1(n169),
	.B0(n488),
	.A1(n328),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U295 (
	.Y(n425),
	.B1(n168),
	.B0(n488),
	.A1(n328),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U296 (
	.Y(n426),
	.B1(n167),
	.B0(n488),
	.A1(n328),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U297 (
	.Y(n427),
	.B1(n166),
	.B0(n488),
	.A1(n328),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U298 (
	.Y(n428),
	.B1(n165),
	.B0(n488),
	.A1(n328),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U299 (
	.Y(n429),
	.B1(n164),
	.B0(n488),
	.A1(n328),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U300 (
	.Y(n430),
	.B1(n163),
	.B0(n488),
	.A1(n328),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U301 (
	.Y(n431),
	.B1(n162),
	.B0(n488),
	.A1(n328),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U302 (
	.Y(n432),
	.B1(n161),
	.B0(n487),
	.A1(n329),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U303 (
	.Y(n433),
	.B1(n160),
	.B0(n487),
	.A1(n329),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U304 (
	.Y(n434),
	.B1(n159),
	.B0(n487),
	.A1(n329),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U305 (
	.Y(n435),
	.B1(n158),
	.B0(n487),
	.A1(n329),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U306 (
	.Y(n436),
	.B1(n157),
	.B0(n487),
	.A1(n329),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U307 (
	.Y(n437),
	.B1(n156),
	.B0(n487),
	.A1(n329),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U308 (
	.Y(n438),
	.B1(n155),
	.B0(n487),
	.A1(n329),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U309 (
	.Y(n439),
	.B1(n154),
	.B0(n487),
	.A1(n329),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U310 (
	.Y(n456),
	.B1(n153),
	.B0(n486),
	.A1(n333),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U311 (
	.Y(n457),
	.B1(n152),
	.B0(n486),
	.A1(n333),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U312 (
	.Y(n458),
	.B1(n151),
	.B0(n486),
	.A1(n333),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U313 (
	.Y(n459),
	.B1(n150),
	.B0(n486),
	.A1(n333),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U314 (
	.Y(n460),
	.B1(n149),
	.B0(n486),
	.A1(n333),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U315 (
	.Y(n461),
	.B1(n148),
	.B0(n486),
	.A1(n333),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U316 (
	.Y(n462),
	.B1(n147),
	.B0(n486),
	.A1(n333),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U317 (
	.Y(n463),
	.B1(n146),
	.B0(n486),
	.A1(n333),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U318 (
	.Y(n464),
	.B1(n145),
	.B0(n485),
	.A1(n334),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U319 (
	.Y(n465),
	.B1(n144),
	.B0(n485),
	.A1(n334),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U320 (
	.Y(n466),
	.B1(n143),
	.B0(n485),
	.A1(n334),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U321 (
	.Y(n467),
	.B1(n142),
	.B0(n485),
	.A1(n334),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U322 (
	.Y(n468),
	.B1(n141),
	.B0(n485),
	.A1(n334),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U323 (
	.Y(n469),
	.B1(n140),
	.B0(n485),
	.A1(n334),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U324 (
	.Y(n470),
	.B1(n139),
	.B0(n485),
	.A1(n334),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U325 (
	.Y(n471),
	.B1(n138),
	.B0(n485),
	.A1(n334),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U326 (
	.Y(n344),
	.B1(n201),
	.B0(n491),
	.A1(n499),
	.A0(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U327 (
	.Y(n345),
	.B1(n200),
	.B0(n491),
	.A1(n500),
	.A0(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U328 (
	.Y(n346),
	.B1(n199),
	.B0(n491),
	.A1(n501),
	.A0(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U329 (
	.Y(n347),
	.B1(n198),
	.B0(n491),
	.A1(n502),
	.A0(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U330 (
	.Y(n348),
	.B1(n197),
	.B0(n491),
	.A1(n503),
	.A0(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U331 (
	.Y(n376),
	.B1(n185),
	.B0(n490),
	.A1(n320),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U332 (
	.Y(n377),
	.B1(n184),
	.B0(n490),
	.A1(n320),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U333 (
	.Y(n378),
	.B1(n183),
	.B0(n490),
	.A1(n320),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U334 (
	.Y(n379),
	.B1(n182),
	.B0(n490),
	.A1(n320),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U335 (
	.Y(n380),
	.B1(n181),
	.B0(n490),
	.A1(n320),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U336 (
	.Y(n381),
	.B1(n180),
	.B0(n490),
	.A1(n320),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U337 (
	.Y(n382),
	.B1(n179),
	.B0(n490),
	.A1(n320),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U338 (
	.Y(n383),
	.B1(n178),
	.B0(n490),
	.A1(n320),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U339 (
	.Y(n384),
	.B1(n177),
	.B0(n489),
	.A1(n322),
	.A0(n499), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U340 (
	.Y(n385),
	.B1(n176),
	.B0(n489),
	.A1(n322),
	.A0(n500), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U341 (
	.Y(n386),
	.B1(n175),
	.B0(n489),
	.A1(n322),
	.A0(n501), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U342 (
	.Y(n387),
	.B1(n174),
	.B0(n489),
	.A1(n322),
	.A0(n502), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U343 (
	.Y(n388),
	.B1(n173),
	.B0(n489),
	.A1(n322),
	.A0(n503), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U344 (
	.Y(n389),
	.B1(n172),
	.B0(n489),
	.A1(n322),
	.A0(n504), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U345 (
	.Y(n390),
	.B1(n171),
	.B0(n489),
	.A1(n322),
	.A0(n505), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U346 (
	.Y(n391),
	.B1(n170),
	.B0(n489),
	.A1(n322),
	.A0(n506), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U347 (
	.Y(n392),
	.B1(n323),
	.B0(n499),
	.A1N(\Reg_File[6][0] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U348 (
	.Y(n393),
	.B1(n323),
	.B0(n500),
	.A1N(\Reg_File[6][1] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U349 (
	.Y(n394),
	.B1(n323),
	.B0(n501),
	.A1N(\Reg_File[6][2] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U350 (
	.Y(n395),
	.B1(n323),
	.B0(n502),
	.A1N(\Reg_File[6][3] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U351 (
	.Y(n396),
	.B1(n323),
	.B0(n503),
	.A1N(\Reg_File[6][4] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U352 (
	.Y(n397),
	.B1(n323),
	.B0(n504),
	.A1N(\Reg_File[6][5] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U353 (
	.Y(n398),
	.B1(n323),
	.B0(n505),
	.A1N(\Reg_File[6][6] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U354 (
	.Y(n399),
	.B1(n323),
	.B0(n506),
	.A1N(\Reg_File[6][7] ),
	.A0N(n323), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U355 (
	.Y(n400),
	.B1(n324),
	.B0(n499),
	.A1N(\Reg_File[7][0] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U356 (
	.Y(n401),
	.B1(n324),
	.B0(n500),
	.A1N(\Reg_File[7][1] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U357 (
	.Y(n402),
	.B1(n324),
	.B0(n501),
	.A1N(\Reg_File[7][2] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U358 (
	.Y(n403),
	.B1(n324),
	.B0(n502),
	.A1N(\Reg_File[7][3] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U359 (
	.Y(n404),
	.B1(n324),
	.B0(n503),
	.A1N(\Reg_File[7][4] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U360 (
	.Y(n405),
	.B1(n324),
	.B0(n504),
	.A1N(\Reg_File[7][5] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U361 (
	.Y(n406),
	.B1(n324),
	.B0(n505),
	.A1N(\Reg_File[7][6] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U362 (
	.Y(n407),
	.B1(n324),
	.B0(n506),
	.A1N(\Reg_File[7][7] ),
	.A0N(n324), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U363 (
	.Y(n361),
	.B1(n318),
	.B0(n500),
	.A1N(REG2[1]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U364 (
	.Y(n362),
	.B1(n318),
	.B0(n501),
	.A1N(REG2[2]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U365 (
	.Y(n363),
	.B1(n318),
	.B0(n502),
	.A1N(REG2[3]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U366 (
	.Y(n364),
	.B1(n318),
	.B0(n503),
	.A1N(REG2[4]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U367 (
	.Y(n366),
	.B1(n318),
	.B0(n505),
	.A1N(REG2[6]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U368 (
	.Y(n367),
	.B1(n318),
	.B0(n506),
	.A1N(REG2[7]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U369 (
	.Y(n368),
	.B1(n319),
	.B0(n499),
	.A1N(REG3[0]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U370 (
	.Y(n369),
	.B1(n319),
	.B0(n500),
	.A1N(REG3[1]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U371 (
	.Y(n370),
	.B1(n319),
	.B0(n501),
	.A1N(REG3[2]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U372 (
	.Y(n371),
	.B1(n319),
	.B0(n502),
	.A1N(REG3[3]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U373 (
	.Y(n372),
	.B1(n319),
	.B0(n503),
	.A1N(REG3[4]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U374 (
	.Y(n374),
	.B1(n319),
	.B0(n505),
	.A1N(REG3[6]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U375 (
	.Y(n375),
	.B1(n319),
	.B0(n506),
	.A1N(REG3[7]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U376 (
	.Y(n408),
	.B1(n325),
	.B0(n499),
	.A1N(\Reg_File[8][0] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U377 (
	.Y(n409),
	.B1(n325),
	.B0(n500),
	.A1N(\Reg_File[8][1] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U378 (
	.Y(n410),
	.B1(n325),
	.B0(n501),
	.A1N(\Reg_File[8][2] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U379 (
	.Y(n411),
	.B1(n325),
	.B0(n502),
	.A1N(\Reg_File[8][3] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U380 (
	.Y(n412),
	.B1(n325),
	.B0(n503),
	.A1N(\Reg_File[8][4] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U381 (
	.Y(n413),
	.B1(n325),
	.B0(n504),
	.A1N(\Reg_File[8][5] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U382 (
	.Y(n414),
	.B1(n325),
	.B0(n505),
	.A1N(\Reg_File[8][6] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U383 (
	.Y(n415),
	.B1(n325),
	.B0(n506),
	.A1N(\Reg_File[8][7] ),
	.A0N(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U384 (
	.Y(n416),
	.B1(n327),
	.B0(n499),
	.A1N(\Reg_File[9][0] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U385 (
	.Y(n417),
	.B1(n327),
	.B0(n500),
	.A1N(\Reg_File[9][1] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U386 (
	.Y(n418),
	.B1(n327),
	.B0(n501),
	.A1N(\Reg_File[9][2] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U387 (
	.Y(n419),
	.B1(n327),
	.B0(n502),
	.A1N(\Reg_File[9][3] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U388 (
	.Y(n420),
	.B1(n327),
	.B0(n503),
	.A1N(\Reg_File[9][4] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U389 (
	.Y(n421),
	.B1(n327),
	.B0(n504),
	.A1N(\Reg_File[9][5] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U390 (
	.Y(n422),
	.B1(n327),
	.B0(n505),
	.A1N(\Reg_File[9][6] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U391 (
	.Y(n423),
	.B1(n327),
	.B0(n506),
	.A1N(\Reg_File[9][7] ),
	.A0N(n327), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U392 (
	.Y(n440),
	.B1(n330),
	.B0(n499),
	.A1N(\Reg_File[12][0] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U393 (
	.Y(n441),
	.B1(n330),
	.B0(n500),
	.A1N(\Reg_File[12][1] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U394 (
	.Y(n442),
	.B1(n330),
	.B0(n501),
	.A1N(\Reg_File[12][2] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U395 (
	.Y(n443),
	.B1(n330),
	.B0(n502),
	.A1N(\Reg_File[12][3] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U396 (
	.Y(n444),
	.B1(n330),
	.B0(n503),
	.A1N(\Reg_File[12][4] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U397 (
	.Y(n445),
	.B1(n330),
	.B0(n504),
	.A1N(\Reg_File[12][5] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U398 (
	.Y(n446),
	.B1(n330),
	.B0(n505),
	.A1N(\Reg_File[12][6] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U399 (
	.Y(n447),
	.B1(n330),
	.B0(n506),
	.A1N(\Reg_File[12][7] ),
	.A0N(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U400 (
	.Y(n448),
	.B1(n332),
	.B0(n499),
	.A1N(\Reg_File[13][0] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U401 (
	.Y(n449),
	.B1(n332),
	.B0(n500),
	.A1N(\Reg_File[13][1] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U402 (
	.Y(n450),
	.B1(n332),
	.B0(n501),
	.A1N(\Reg_File[13][2] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U403 (
	.Y(n451),
	.B1(n332),
	.B0(n502),
	.A1N(\Reg_File[13][3] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U404 (
	.Y(n452),
	.B1(n332),
	.B0(n503),
	.A1N(\Reg_File[13][4] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U405 (
	.Y(n453),
	.B1(n332),
	.B0(n504),
	.A1N(\Reg_File[13][5] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U406 (
	.Y(n454),
	.B1(n332),
	.B0(n505),
	.A1N(\Reg_File[13][6] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U407 (
	.Y(n455),
	.B1(n332),
	.B0(n506),
	.A1N(\Reg_File[13][7] ),
	.A0N(n332), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U408 (
	.Y(n360),
	.B1(n318),
	.B0(n499),
	.A1N(REG2[0]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U409 (
	.Y(n365),
	.B1(n318),
	.B0(n504),
	.A1N(REG2[5]),
	.A0N(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U410 (
	.Y(n373),
	.B1(n319),
	.B0(n504),
	.A1N(REG3[5]),
	.A0N(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U411 (
	.Y(n353),
	.S0(n186),
	.B(WrData[1]),
	.A(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U412 (
	.Y(n483),
	.B1(n495),
	.B0(REG3[0]),
	.A1(n493),
	.A0(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U413 (
	.Y(n482),
	.B1(n495),
	.B0(REG3[1]),
	.A1(n493),
	.A0(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U414 (
	.Y(n480),
	.B1(n495),
	.B0(REG3[2]),
	.A1(n493),
	.A0(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U415 (
	.Y(n478),
	.B1(n495),
	.B0(REG3[3]),
	.A1(n493),
	.A0(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U416 (
	.Y(n476),
	.B1(n495),
	.B0(REG3[4]),
	.A1(n493),
	.A0(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U417 (
	.Y(n473),
	.B1(n495),
	.B0(REG3[5]),
	.A1(n493),
	.A0(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U418 (
	.Y(n310),
	.B1(n495),
	.B0(REG3[6]),
	.A1(n493),
	.A0(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U419 (
	.Y(n290),
	.B1(n495),
	.B0(REG3[7]),
	.A1(n493),
	.A0(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U420 (
	.Y(n240),
	.B1(n242),
	.B0(\Reg_File[13][0] ),
	.A1(n241),
	.A0(\Reg_File[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U421 (
	.Y(n243),
	.B1(n242),
	.B0(\Reg_File[9][0] ),
	.A1(n241),
	.A0(\Reg_File[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U422 (
	.Y(n252),
	.B1(n242),
	.B0(\Reg_File[13][1] ),
	.A1(n241),
	.A0(\Reg_File[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U423 (
	.Y(n253),
	.B1(n242),
	.B0(\Reg_File[9][1] ),
	.A1(n241),
	.A0(\Reg_File[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U424 (
	.Y(n262),
	.B1(n242),
	.B0(\Reg_File[13][2] ),
	.A1(n241),
	.A0(\Reg_File[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U425 (
	.Y(n263),
	.B1(n242),
	.B0(\Reg_File[9][2] ),
	.A1(n241),
	.A0(\Reg_File[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U426 (
	.Y(n272),
	.B1(n242),
	.B0(\Reg_File[13][3] ),
	.A1(n241),
	.A0(\Reg_File[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U427 (
	.Y(n273),
	.B1(n242),
	.B0(\Reg_File[9][3] ),
	.A1(n241),
	.A0(\Reg_File[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U428 (
	.Y(n282),
	.B1(n242),
	.B0(\Reg_File[13][4] ),
	.A1(n241),
	.A0(\Reg_File[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U429 (
	.Y(n283),
	.B1(n242),
	.B0(\Reg_File[9][4] ),
	.A1(n241),
	.A0(\Reg_File[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U430 (
	.Y(n292),
	.B1(n242),
	.B0(\Reg_File[13][5] ),
	.A1(n241),
	.A0(\Reg_File[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U431 (
	.Y(n293),
	.B1(n242),
	.B0(\Reg_File[9][5] ),
	.A1(n241),
	.A0(\Reg_File[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U432 (
	.Y(n302),
	.B1(n242),
	.B0(\Reg_File[13][6] ),
	.A1(n241),
	.A0(\Reg_File[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U433 (
	.Y(n303),
	.B1(n242),
	.B0(\Reg_File[9][6] ),
	.A1(n241),
	.A0(\Reg_File[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U434 (
	.Y(n312),
	.B1(n242),
	.B0(\Reg_File[13][7] ),
	.A1(n241),
	.A0(\Reg_File[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U435 (
	.Y(n313),
	.B1(n242),
	.B0(\Reg_File[9][7] ),
	.A1(n241),
	.A0(\Reg_File[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U436 (
	.Y(n343),
	.B0(n226),
	.A1N(n314),
	.A0N(RdData_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U437 (
	.Y(REG1[2]),
	.A(n191), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U441 (
	.Y(n309),
	.C0(n290),
	.B1(n242),
	.B0(REG1[7]),
	.A1(n241),
	.A0(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U442 (
	.Y(n359),
	.S0(n186),
	.B(WrData[7]),
	.A(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U443 (
	.Y(n358),
	.S0(n186),
	.B(WrData[6]),
	.A(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U444 (
	.Y(n299),
	.C0(n310),
	.B1(n242),
	.B0(REG1[6]),
	.A1(n241),
	.A0(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U445 (
	.Y(n351),
	.S0(n491),
	.B(WrData[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U446 (
	.Y(n563),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U447 (
	.Y(n564),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U448 (
	.Y(n565),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U449 (
	.Y(n566),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_test_1 (
	A, 
	B, 
	ALU_FUN, 
	EN, 
	CLK, 
	RST, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input EN;
   input CLK;
   input RST;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N157;
   wire N158;
   wire N159;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n53;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n71;
   wire n72;
   wire n73;
   wire n77;
   wire n78;
   wire n79;
   wire n83;
   wire n84;
   wire n85;
   wire n89;
   wire n90;
   wire n91;
   wire n95;
   wire n96;
   wire n97;
   wire n105;
   wire n106;
   wire n107;
   wire n109;
   wire n118;
   wire n120;
   wire n121;
   wire n123;
   wire n3;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n27;
   wire n32;
   wire n33;
   wire n34;
   wire n46;
   wire n47;
   wire n52;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n74;
   wire n75;
   wire n76;
   wire n80;
   wire n81;
   wire n82;
   wire n86;
   wire n87;
   wire n88;
   wire n92;
   wire n93;
   wire n94;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n108;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n119;
   wire n122;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire [15:0] ALU_OUT_Comb;

   // Module instantiations
   CLKINVX2M FE_RC_5_0 (
	.Y(n32),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_RC_4_0 (
	.Y(n33),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[7]),
	.D(ALU_OUT_Comb[7]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[6]),
	.D(ALU_OUT_Comb[6]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[5]),
	.D(ALU_OUT_Comb[5]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[4]),
	.D(ALU_OUT_Comb[4]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[3]),
	.D(ALU_OUT_Comb[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[2]),
	.D(ALU_OUT_Comb[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[15]),
	.D(ALU_OUT_Comb[15]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[14]),
	.D(ALU_OUT_Comb[14]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[13]),
	.D(ALU_OUT_Comb[13]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[12]),
	.D(ALU_OUT_Comb[12]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[11]),
	.D(ALU_OUT_Comb[11]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[10]),
	.D(ALU_OUT_Comb[10]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[9]),
	.D(ALU_OUT_Comb[9]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(ALU_OUT_Comb[8]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[0]),
	.D(ALU_OUT_Comb[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M OUT_VALID_reg (
	.SI(ALU_OUT[15]),
	.SE(test_se),
	.RN(RST),
	.Q(OUT_VALID),
	.D(EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[1]),
	.D(ALU_OUT_Comb[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n144),
	.B1(n27),
	.B0(N92),
	.A1(n148),
	.A0(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U32 (
	.Y(n3),
	.B(n111),
	.A(n120), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n6),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U39 (
	.Y(n8),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U40 (
	.Y(n128),
	.B(n102),
	.A(N125), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n130),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n133),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n150),
	.A(n129), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n142),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n149),
	.A(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n152),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U47 (
	.Y(ALU_OUT_Comb[14]),
	.B0(n49),
	.A1N(n48),
	.A0N(N123), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U48 (
	.Y(ALU_OUT_Comb[13]),
	.B0(n49),
	.A1N(n48),
	.A0N(N122), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U49 (
	.Y(ALU_OUT_Comb[15]),
	.B0(n49),
	.A1N(n48),
	.A0N(N124), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U50 (
	.Y(ALU_OUT_Comb[9]),
	.B0(n49),
	.A1N(n48),
	.A0N(N118), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U51 (
	.Y(ALU_OUT_Comb[10]),
	.B0(n49),
	.A1N(n48),
	.A0N(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U52 (
	.Y(ALU_OUT_Comb[11]),
	.B0(n49),
	.A1N(n48),
	.A0N(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U53 (
	.Y(ALU_OUT_Comb[12]),
	.B0(n49),
	.A1N(n48),
	.A0N(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U54 (
	.Y(n64),
	.B0(n118),
	.A1N(n153),
	.A0N(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U55 (
	.Y(n65),
	.B0(n118),
	.A1N(n154),
	.A0N(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U56 (
	.Y(n129),
	.B(n55),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U57 (
	.Y(n154),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U58 (
	.Y(n116),
	.C(n55),
	.B(n153),
	.AN(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U59 (
	.Y(n135),
	.B(n46),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U60 (
	.Y(n131),
	.B(n129),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U61 (
	.Y(n148),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U62 (
	.Y(n52),
	.C(n55),
	.B(n151),
	.AN(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U63 (
	.Y(n9),
	.B(n47),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U64 (
	.Y(n27),
	.B(n54),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U65 (
	.Y(n54),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U66 (
	.Y(n134),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U67 (
	.Y(n151),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U68 (
	.Y(n153),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U69 (
	.Y(n48),
	.B(n191),
	.AN(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U70 (
	.Y(n88),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U71 (
	.Y(n126),
	.B(n124),
	.A(n125), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U72 (
	.Y(n127),
	.B(n112),
	.A(n113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U73 (
	.Y(ALU_OUT_Comb[7]),
	.B0(n191),
	.A2(n99),
	.A1(n100),
	.A0(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U74 (
	.Y(ALU_OUT_Comb[8]),
	.B0(n191),
	.A1(n51),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U75 (
	.Y(n50),
	.B0(n190),
	.A1(n27),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U76 (
	.Y(n51),
	.B1(n148),
	.B0(N117),
	.A1N(n53),
	.A0N(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U77 (
	.Y(n55),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U78 (
	.Y(n46),
	.B(n55),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U79 (
	.Y(n53),
	.C(n150),
	.B(ALU_FUN[3]),
	.AN(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U80 (
	.Y(n123),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U81 (
	.Y(n140),
	.C(n154),
	.B(ALU_FUN[3]),
	.AN(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U82 (
	.Y(n106),
	.C(n156),
	.B(ALU_FUN[2]),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U83 (
	.Y(n63),
	.C(ALU_FUN[3]),
	.B(n157),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U84 (
	.Y(n49),
	.B(n190),
	.A(EN), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U85 (
	.Y(n190),
	.A(n109), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U86 (
	.Y(n109),
	.C0(n64),
	.B0(n149),
	.A1(n9),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U87 (
	.Y(n157),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U88 (
	.Y(n47),
	.B(n157),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U89 (
	.Y(n56),
	.B(ALU_FUN[3]),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U90 (
	.Y(n156),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U91 (
	.Y(n118),
	.C(ALU_FUN[3]),
	.B(ALU_FUN[0]),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U92 (
	.Y(n107),
	.D(n157),
	.C(ALU_FUN[3]),
	.B(n154),
	.A(N159), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U93 (
	.Y(n74),
	.B1(n149),
	.B0(n197),
	.A1(n27),
	.A0(N95), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U94 (
	.Y(n81),
	.B1(n149),
	.B0(n196),
	.A1(n27),
	.A0(N96), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U95 (
	.Y(n92),
	.B1(n149),
	.B0(n195),
	.A1(n27),
	.A0(N97), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U96 (
	.Y(n121),
	.C(ALU_FUN[0]),
	.B(ALU_FUN[2]),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n191),
	.A(EN), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U98 (
	.Y(n113),
	.A(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U99 (
	.Y(ALU_OUT_Comb[2]),
	.B0(n191),
	.A2(n58),
	.A1(n59),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U100 (
	.Y(n59),
	.B1(A[2]),
	.B0(n152),
	.A1(n9),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U101 (
	.Y(n58),
	.C0(n95),
	.B0(n57),
	.A1(n148),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U102 (
	.Y(n66),
	.B1(n142),
	.B0(N127),
	.A1(n88),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U104 (
	.Y(ALU_OUT_Comb[3]),
	.B0(n191),
	.A2(n68),
	.A1(n69),
	.A0(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U105 (
	.Y(n69),
	.B1(n152),
	.B0(A[3]),
	.A1(n9),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U106 (
	.Y(n68),
	.C0(n89),
	.B0(n67),
	.A1(n148),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U107 (
	.Y(n70),
	.B1(n142),
	.B0(N128),
	.A1(n88),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U108 (
	.Y(ALU_OUT_Comb[4]),
	.B0(n191),
	.A2(n75),
	.A1(n76),
	.A0(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U109 (
	.Y(n76),
	.B1(n152),
	.B0(A[4]),
	.A1(n9),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U110 (
	.Y(n75),
	.C0(n83),
	.B0(n74),
	.A1(n148),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U112 (
	.Y(n94),
	.B1(n152),
	.B0(A[6]),
	.A1(n9),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U113 (
	.Y(n93),
	.C0(n71),
	.B0(n92),
	.A1(n148),
	.A0(N115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U114 (
	.Y(ALU_OUT_Comb[5]),
	.B0(n191),
	.A2(n82),
	.A1(n86),
	.A0(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U115 (
	.Y(n86),
	.B1(n152),
	.B0(A[5]),
	.A1(n9),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U116 (
	.Y(n87),
	.B1(n142),
	.B0(N130),
	.A1(n88),
	.A0(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U117 (
	.Y(n82),
	.C0(n77),
	.B0(n81),
	.A1(n148),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U118 (
	.Y(n187),
	.A(n169), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U119 (
	.Y(n124),
	.C(n119),
	.B(n3),
	.A(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U120 (
	.Y(n112),
	.B(n3),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U121 (
	.Y(n72),
	.C0(n152),
	.B1(n65),
	.B0(A[6]),
	.A1(n195),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U122 (
	.Y(n73),
	.C0(n149),
	.B1(n195),
	.B0(n64),
	.A1(n63),
	.A0(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U123 (
	.Y(n83),
	.C1(n198),
	.C0(n53),
	.B1(n85),
	.B0(n34),
	.A1(n32),
	.A0(n84), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U124 (
	.Y(n85),
	.C0(n149),
	.B1(n197),
	.B0(n64),
	.A1(n63),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U125 (
	.Y(n84),
	.C0(n152),
	.B1(n65),
	.B0(A[4]),
	.A1(n197),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U126 (
	.Y(n77),
	.C1(n197),
	.C0(n53),
	.B1(n79),
	.B0(B[5]),
	.A1(n193),
	.A0(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U127 (
	.Y(n193),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U128 (
	.Y(n79),
	.C0(n149),
	.B1(n196),
	.B0(n64),
	.A1(n63),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U129 (
	.Y(n78),
	.C0(n152),
	.B1(n65),
	.B0(A[5]),
	.A1(n196),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U130 (
	.Y(n125),
	.D(n114),
	.C(n115),
	.B(n116),
	.A(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U131 (
	.Y(n102),
	.C(n117),
	.B(n119),
	.A(n115), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U132 (
	.Y(n114),
	.B(n140),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U133 (
	.Y(n143),
	.S0(B[1]),
	.B(n152),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U134 (
	.Y(n132),
	.S0(B[1]),
	.B(n134),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U135 (
	.Y(n137),
	.B(n135),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U136 (
	.Y(n136),
	.S0(B[1]),
	.B(n133),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U137 (
	.Y(n57),
	.B1(n149),
	.B0(n199),
	.A1(n27),
	.A0(N93), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U138 (
	.Y(n67),
	.B1(n149),
	.B0(n198),
	.A1(n27),
	.A0(N94), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U140 (
	.Y(n122),
	.B(n148),
	.A(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U141 (
	.Y(n197),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U142 (
	.Y(n198),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U143 (
	.Y(n199),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U144 (
	.Y(n195),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U145 (
	.Y(n196),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U146 (
	.Y(ALU_OUT_Comb[1]),
	.B0(n191),
	.A1(n146),
	.A0(n147), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U147 (
	.Y(n146),
	.C0(n143),
	.B0(n144),
	.A1(n145),
	.A0(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U148 (
	.Y(n145),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U152 (
	.Y(n141),
	.C0(n139),
	.B0(n105),
	.A1N(A[2]),
	.A0(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U153 (
	.Y(n139),
	.S0(A[1]),
	.B(n137),
	.A(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U154 (
	.Y(n105),
	.B0(n107),
	.A2(n106),
	.A1(ALU_FUN[3]),
	.A0(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U155 (
	.Y(n138),
	.B(n131),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U156 (
	.Y(n155),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U157 (
	.Y(n111),
	.S0(A[0]),
	.B(n108),
	.A(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U158 (
	.Y(n120),
	.B0(n107),
	.A2(n121),
	.A1(ALU_FUN[3]),
	.A0(N157), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U159 (
	.Y(n110),
	.B(n131),
	.A(n103), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U160 (
	.Y(n108),
	.B(n135),
	.A(n104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U161 (
	.Y(n96),
	.C0(n152),
	.B1(n65),
	.B0(A[2]),
	.A1(n199),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U162 (
	.Y(n97),
	.C0(n149),
	.B1(n199),
	.B0(n64),
	.A1(n63),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U163 (
	.Y(n90),
	.C0(n152),
	.B1(n65),
	.B0(A[3]),
	.A1(n198),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U164 (
	.Y(n91),
	.C0(n149),
	.B1(n198),
	.B0(n64),
	.A1(n63),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U165 (
	.Y(n185),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n115),
	.B(n9),
	.A(N100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n119),
	.B(n27),
	.A(N91), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21XLM U168 (
	.Y(n159),
	.B0(B[1]),
	.A1(n155),
	.A0(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U169 (
	.Y(n188),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U170 (
	.Y(ALU_OUT_Comb[0]),
	.C0(n191),
	.B0(n126),
	.A1(n127),
	.A0(n128), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222XLM U171 (
	.Y(n95),
	.C1(n155),
	.C0(n53),
	.B1(n97),
	.B0(n8),
	.A1(n186),
	.A0(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U172 (
	.Y(n186),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U173 (
	.Y(n194),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U174 (
	.Y(ALU_OUT_Comb[6]),
	.B0(n191),
	.A2(n93),
	.A1(n94),
	.A0(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U175 (
	.Y(n100),
	.B1(A[7]),
	.B0(n131),
	.A1(n194),
	.A0(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U176 (
	.Y(n101),
	.B1(n9),
	.B0(N107),
	.A1(n142),
	.A0(N132), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U177 (
	.Y(n99),
	.C0(n60),
	.B1(n148),
	.B0(N116),
	.A1(n27),
	.A0(N98), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U178 (
	.Y(n189),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U179 (
	.Y(n192),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222XLM U180 (
	.Y(n71),
	.C1(n196),
	.C0(n53),
	.B1(n73),
	.B0(B[6]),
	.A1(n189),
	.A0(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32XLM U181 (
	.Y(n165),
	.B1(n195),
	.B0(B[6]),
	.A2(n177),
	.A1(n174),
	.A0(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2XLM U182 (
	.Y(n177),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U183 (
	.Y(n34),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U184 (
	.Y(n98),
	.B1(n142),
	.B0(N131),
	.A1(n88),
	.A0(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U185 (
	.Y(n61),
	.C0(n152),
	.B1(n65),
	.B0(A[7]),
	.A1(n194),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U186 (
	.Y(n62),
	.C0(n149),
	.B1(n194),
	.B0(n64),
	.A1(A[7]),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222XLM U187 (
	.Y(n89),
	.C1(n199),
	.C0(n53),
	.B1(n91),
	.B0(B[3]),
	.A1(n188),
	.A0(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U188 (
	.Y(n181),
	.B(n194),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U189 (
	.Y(n104),
	.S0(B[0]),
	.B(n133),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U190 (
	.Y(n117),
	.S0(B[0]),
	.B(n135),
	.A(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U191 (
	.Y(n103),
	.S0(B[0]),
	.B(n134),
	.A(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U192 (
	.Y(n184),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222XLM U193 (
	.Y(n60),
	.C1(n195),
	.C0(n53),
	.B1(n62),
	.B0(B[7]),
	.A1(n192),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U194 (
	.Y(n180),
	.B(B[7]),
	.A(n194), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U195 (
	.Y(n147),
	.C0(n141),
	.B1(n9),
	.B0(N101),
	.A1(n142),
	.A0(N126), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22XLM U196 (
	.Y(n80),
	.B1(n142),
	.B0(N129),
	.A1(n88),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U197 (
	.Y(n173),
	.B(A[4]),
	.AN(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U198 (
	.Y(n162),
	.B(n34),
	.AN(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U199 (
	.Y(n175),
	.B(n162),
	.A(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U200 (
	.Y(n170),
	.B(A[3]),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U201 (
	.Y(n161),
	.B(A[2]),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U202 (
	.Y(n158),
	.B(A[0]),
	.A(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U203 (
	.Y(n172),
	.B(n186),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U204 (
	.Y(n167),
	.B(n172),
	.AN(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U205 (
	.Y(n160),
	.C0(n159),
	.B0(n167),
	.A1(n185),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U206 (
	.Y(n171),
	.B(n188),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U207 (
	.Y(n163),
	.B0(n171),
	.A2(n160),
	.A1(n161),
	.A0(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U208 (
	.Y(n178),
	.B(B[5]),
	.AN(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U209 (
	.Y(n164),
	.C0(n178),
	.B0(n162),
	.A1(n163),
	.A0(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U210 (
	.Y(n174),
	.B(A[5]),
	.AN(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U211 (
	.Y(N159),
	.B0(n181),
	.A1(n165),
	.A0(n180), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U212 (
	.Y(n168),
	.B(n184),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U213 (
	.Y(n166),
	.B0(B[1]),
	.A1(n155),
	.A0(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U214 (
	.Y(n169),
	.C0(n166),
	.B0(n167),
	.A1(n155),
	.A0(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U215 (
	.Y(n176),
	.B0(n170),
	.A2(n171),
	.A1(n172),
	.A0(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U216 (
	.Y(n179),
	.C0(n173),
	.B0(n174),
	.A1N(n176),
	.A0(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U217 (
	.Y(n182),
	.B1(n189),
	.B0(A[6]),
	.A2(n177),
	.A1(n178),
	.A0(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U218 (
	.Y(n183),
	.B0(n180),
	.A1N(n182),
	.A0(n181), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U219 (
	.Y(N158),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U220 (
	.Y(N157),
	.B(N158),
	.A(N159), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_sub_0 sub_52 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		n34,
		B[3],
		n8,
		B[1],
		B[0] }),
	.CI(1'b0),
	.DIFF({ N108,
		N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100 }),
	.n184(n184),
	.n189(n189),
	.n188(n188),
	.n193(n193),
	.n186(n186),
	.n192(n192), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_0 add_48 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		n34,
		B[3],
		n8,
		B[1],
		B[0] }),
	.CI(1'b0),
	.SUM({ N99,
		N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW02_mult_0 mult_56 (
	.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ B[7],
		B[6],
		B[5],
		n34,
		B[3],
		n8,
		B[1],
		B[0] }),
	.TC(1'b0),
	.PRODUCT({ N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109 }),
	.n196(n196),
	.n195(n195),
	.n155(n155),
	.n199(n199),
	.n198(n198),
	.n197(n197),
	.n193(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW_div_uns_1 div_60 (
	.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.b({ B[7],
		B[6],
		B[5],
		n33,
		B[3],
		n7,
		B[1],
		B[0] }),
	.quotient({ N132,
		N131,
		N130,
		N129,
		N128,
		N127,
		N126,
		N125 }),
	.n196(n196),
	.n155(n155),
	.n199(n199),
	.n197(n197),
	.n193(n193), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n184, 
	n189, 
	n188, 
	n193, 
	n186, 
	n192, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n184;
   input n189;
   input n188;
   input n193;
   input n186;
   input n192;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n5;
   wire n8;
   wire [9:0] carry;

   // Module instantiations
   ADDFXLM U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n192),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n8),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n188),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n186),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n189),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n193),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n5),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(n5),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(carry[1]),
	.B(n1),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n1),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U6 (
	.Y(n8),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire [8:1] carry;

   // Module instantiations
   ADDFX1M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2XLM U2 (
	.Y(SUM[0]),
	.B(n2),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n2),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n196, 
	n195, 
	n155, 
	n199, 
	n198, 
	n197, 
	n193, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n196;
   input n195;
   input n155;
   input n199;
   input n198;
   input n197;
   input n193;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   // Module instantiations
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n7),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n4),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n9),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n6),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n5),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n8),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n3),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U10 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U11 (
	.Y(n11),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n27),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U14 (
	.Y(n12),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n23),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n22),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n20),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n19),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n18),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n21),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U26 (
	.Y(\SUMB[1][2] ),
	.B(n19),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U27 (
	.Y(\SUMB[1][6] ),
	.B(n23),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U28 (
	.Y(\SUMB[1][5] ),
	.B(n22),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n13),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U30 (
	.Y(n14),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U31 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U34 (
	.Y(n16),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][4] ),
	.B(n21),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U36 (
	.Y(\SUMB[1][3] ),
	.B(n20),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U37 (
	.Y(\SUMB[1][1] ),
	.B(n18),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n37),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n35),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n36),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n39),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n38),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U46 (
	.Y(n30),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U47 (
	.Y(n28),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U48 (
	.Y(n29),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U49 (
	.Y(n32),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n25),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U51 (
	.Y(n31),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U52 (
	.Y(n24),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(\ab[7][7] ),
	.B(n24),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][6] ),
	.B(n25),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][5] ),
	.B(n193),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][4] ),
	.B(n27),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][3] ),
	.B(n28),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][2] ),
	.B(n29),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][1] ),
	.B(n30),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][0] ),
	.B(n31),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[6][7] ),
	.B(n195),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][6] ),
	.B(n195),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][5] ),
	.B(n195),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][4] ),
	.B(n195),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][3] ),
	.B(n195),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][2] ),
	.B(n195),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][1] ),
	.B(n195),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][0] ),
	.B(n195),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[5][7] ),
	.B(n196),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][6] ),
	.B(n196),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][5] ),
	.B(n196),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][4] ),
	.B(n196),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][3] ),
	.B(n196),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][2] ),
	.B(n196),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][1] ),
	.B(n196),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][0] ),
	.B(n196),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[4][7] ),
	.B(n35),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][6] ),
	.B(n35),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][5] ),
	.B(n35),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][4] ),
	.B(n35),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][3] ),
	.B(n35),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][2] ),
	.B(n35),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][1] ),
	.B(n35),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][0] ),
	.B(n35),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[3][7] ),
	.B(n36),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][6] ),
	.B(n36),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][5] ),
	.B(n36),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][4] ),
	.B(n36),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][3] ),
	.B(n36),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][2] ),
	.B(n36),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][1] ),
	.B(n36),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][0] ),
	.B(n36),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[2][7] ),
	.B(n37),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][6] ),
	.B(n37),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][5] ),
	.B(n37),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][4] ),
	.B(n37),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][3] ),
	.B(n37),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][2] ),
	.B(n37),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][1] ),
	.B(n37),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][0] ),
	.B(n37),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[1][7] ),
	.B(n38),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][6] ),
	.B(n38),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][5] ),
	.B(n38),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][4] ),
	.B(n38),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][3] ),
	.B(n38),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][2] ),
	.B(n38),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][1] ),
	.B(n38),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][0] ),
	.B(n38),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[0][7] ),
	.B(n39),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][6] ),
	.B(n39),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][5] ),
	.B(n39),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][4] ),
	.B(n39),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][3] ),
	.B(n39),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][2] ),
	.B(n39),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][1] ),
	.B(n39),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(PRODUCT[0]),
	.B(n39),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n12,
		n11,
		n16,
		n15,
		n14,
		n13,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n19),
	.A1(A[12]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n15),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(SUM[7]),
	.B(n8),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n8),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(SUM[6]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n9),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U9 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U10 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U12 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U13 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(SUM[9]),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(SUM[8]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U18 (
	.Y(n14),
	.B(n17),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n19),
	.B0(B[12]),
	.A1(n18),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U20 (
	.Y(SUM[12]),
	.C(n18),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U21 (
	.Y(n18),
	.B0N(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U22 (
	.Y(SUM[11]),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n20),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U25 (
	.Y(n22),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U26 (
	.Y(n21),
	.B0(n26),
	.A1(n25),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(SUM[10]),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U28 (
	.Y(n25),
	.B0(n12),
	.A1N(n13),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U29 (
	.Y(n12),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(n13),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U31 (
	.Y(n10),
	.B0(n17),
	.A1(n16),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n17),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(n16),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n27),
	.B(n26),
	.AN(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n26),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U36 (
	.Y(n24),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW_div_uns_1 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n196, 
	n155, 
	n199, 
	n197, 
	n193, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n196;
   input n155;
   input n199;
   input n197;
   input n193;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire FE_RN_665_0;
   wire FE_RN_663_0;
   wire FE_RN_662_0;
   wire FE_RN_661_0;
   wire FE_RN_660_0;
   wire FE_RN_659_0;
   wire FE_RN_658_0;
   wire FE_RN_657_0;
   wire FE_RN_656_0;
   wire FE_RN_655_0;
   wire FE_RN_654_0;
   wire FE_RN_652_0;
   wire FE_RN_651_0;
   wire FE_RN_650_0;
   wire FE_RN_649_0;
   wire FE_RN_648_0;
   wire FE_RN_647_0;
   wire FE_RN_646_0;
   wire FE_RN_645_0;
   wire FE_RN_644_0;
   wire FE_RN_643_0;
   wire FE_RN_641_0;
   wire FE_RN_640_0;
   wire FE_RN_639_0;
   wire FE_RN_638_0;
   wire FE_RN_636_0;
   wire FE_RN_635_0;
   wire FE_RN_633_0;
   wire FE_RN_632_0;
   wire FE_RN_631_0;
   wire FE_RN_630_0;
   wire FE_RN_629_0;
   wire FE_RN_603_0;
   wire FE_RN_602_0;
   wire FE_RN_601_0;
   wire FE_RN_600_0;
   wire FE_RN_599_0;
   wire FE_RN_598_0;
   wire FE_RN_597_0;
   wire FE_RN_596_0;
   wire FE_RN_595_0;
   wire FE_RN_592_0;
   wire FE_RN_591_0;
   wire FE_RN_590_0;
   wire FE_RN_589_0;
   wire FE_RN_588_0;
   wire FE_RN_587_0;
   wire FE_RN_586_0;
   wire FE_RN_585_0;
   wire FE_RN_584_0;
   wire FE_RN_583_0;
   wire FE_RN_582_0;
   wire FE_RN_581_0;
   wire FE_RN_580_0;
   wire FE_RN_579_0;
   wire FE_RN_578_0;
   wire FE_RN_576_0;
   wire FE_RN_575_0;
   wire FE_RN_574_0;
   wire FE_RN_573_0;
   wire FE_RN_572_0;
   wire FE_RN_571_0;
   wire FE_RN_570_0;
   wire FE_RN_568_0;
   wire FE_RN_566_0;
   wire FE_RN_565_0;
   wire FE_RN_564_0;
   wire FE_RN_563_0;
   wire FE_RN_562_0;
   wire FE_RN_541_0;
   wire FE_RN_540_0;
   wire FE_RN_528_0;
   wire FE_RN_527_0;
   wire FE_RN_526_0;
   wire FE_RN_525_0;
   wire FE_RN_523_0;
   wire FE_RN_522_0;
   wire FE_RN_521_0;
   wire FE_RN_520_0;
   wire FE_RN_519_0;
   wire FE_RN_518_0;
   wire FE_RN_516_0;
   wire FE_RN_515_0;
   wire FE_RN_514_0;
   wire FE_RN_513_0;
   wire FE_RN_512_0;
   wire FE_RN_511_0;
   wire FE_RN_509_0;
   wire FE_RN_508_0;
   wire FE_RN_507_0;
   wire FE_RN_506_0;
   wire FE_RN_505_0;
   wire FE_RN_503_0;
   wire FE_RN_502_0;
   wire FE_RN_501_0;
   wire FE_RN_500_0;
   wire FE_RN_499_0;
   wire FE_RN_498_0;
   wire FE_RN_497_0;
   wire FE_RN_495_0;
   wire FE_RN_493_0;
   wire FE_RN_492_0;
   wire FE_RN_491_0;
   wire FE_RN_490_0;
   wire FE_RN_147_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_59_0;
   wire FE_RN_58_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_RN_47_0;
   wire FE_RN_45_0;
   wire FE_RN_44_0;
   wire FE_RN_43_0;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_33_0;
   wire FE_RN_32_0;
   wire FE_RN_31_0;
   wire FE_OFN11_u_div_BInv_2_;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[6][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n24;
   wire n26;
   wire n28;
   wire n29;
   wire n31;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n45;
   wire n48;
   wire n49;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire [7:0] \u_div/BInv ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_819_0 (
	.Y(FE_RN_665_0),
	.A(FE_RN_656_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_817_0 (
	.Y(FE_RN_663_0),
	.A(FE_RN_638_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_816_0 (
	.Y(FE_RN_662_0),
	.B0(FE_RN_640_0),
	.A1(FE_RN_635_0),
	.A0(FE_RN_663_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_815_0 (
	.Y(FE_RN_661_0),
	.B0(FE_RN_662_0),
	.A1N(FE_RN_635_0),
	.A0N(FE_RN_630_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_814_0 (
	.Y(FE_RN_660_0),
	.B(FE_RN_665_0),
	.A(FE_RN_661_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_813_0 (
	.Y(FE_RN_659_0),
	.A(FE_RN_644_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_812_0 (
	.Y(FE_RN_658_0),
	.B(FE_RN_659_0),
	.A(FE_RN_650_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_811_0 (
	.Y(FE_RN_657_0),
	.A(FE_RN_635_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M FE_RC_810_0 (
	.Y(FE_RN_656_0),
	.B(\u_div/BInv [6]),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_809_0 (
	.Y(FE_RN_655_0),
	.B0(FE_RN_656_0),
	.A1(FE_RN_657_0),
	.A0(FE_RN_658_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_808_0 (
	.Y(\u_div/SumTmp[1][6] ),
	.B(FE_RN_660_0),
	.A(FE_RN_655_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_807_0 (
	.Y(FE_RN_654_0),
	.B(\u_div/BInv [5]),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_805_0 (
	.Y(FE_RN_652_0),
	.B(FE_RN_659_0),
	.AN(FE_RN_635_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_804_0 (
	.Y(FE_RN_651_0),
	.B(FE_RN_643_0),
	.A(FE_RN_638_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_803_0 (
	.Y(FE_RN_650_0),
	.B(FE_RN_586_0),
	.A(FE_RN_651_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_802_0 (
	.Y(\u_div/SumTmp[1][5] ),
	.S0(FE_RN_650_0),
	.B(FE_RN_652_0),
	.A(FE_RN_654_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_801_0 (
	.Y(FE_RN_649_0),
	.A(\u_div/BInv [6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_800_0 (
	.Y(FE_RN_648_0),
	.A(FE_RN_643_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_799_0 (
	.Y(FE_RN_647_0),
	.B(FE_RN_648_0),
	.A(FE_RN_635_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_798_0 (
	.Y(FE_RN_646_0),
	.C(FE_RN_649_0),
	.B(FE_RN_644_0),
	.A(FE_RN_647_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_797_0 (
	.Y(FE_RN_645_0),
	.B(\u_div/PartRem[2][6] ),
	.A(FE_RN_646_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_796_0 (
	.Y(FE_RN_644_0),
	.B(\u_div/BInv [5]),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_795_0 (
	.Y(FE_RN_643_0),
	.B(\u_div/BInv [4]),
	.A(FE_RN_595_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_793_0 (
	.Y(FE_RN_641_0),
	.B(FE_RN_648_0),
	.A(FE_RN_635_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_792_0 (
	.Y(FE_RN_640_0),
	.B(FE_RN_644_0),
	.A(FE_RN_641_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_791_0 (
	.Y(FE_RN_639_0),
	.B(\u_div/BInv [6]),
	.A(FE_RN_640_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_790_0 (
	.Y(FE_RN_638_0),
	.B(\u_div/PartRem[2][4] ),
	.A(FE_RN_596_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_788_0 (
	.Y(FE_RN_636_0),
	.A(\u_div/BInv [5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_787_0 (
	.Y(FE_RN_635_0),
	.B(FE_RN_636_0),
	.AN(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_785_0 (
	.Y(FE_RN_633_0),
	.B(FE_RN_649_0),
	.AN(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_784_0 (
	.Y(FE_RN_632_0),
	.A(FE_RN_633_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_783_0 (
	.Y(FE_RN_631_0),
	.B(FE_RN_632_0),
	.AN(FE_RN_635_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_782_0 (
	.Y(FE_RN_630_0),
	.A(FE_RN_586_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X2M FE_RC_781_0 (
	.Y(FE_RN_629_0),
	.B1(FE_RN_630_0),
	.B0(FE_RN_631_0),
	.A2(FE_RN_633_0),
	.A1(FE_RN_635_0),
	.A0(FE_RN_663_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_780_0 (
	.Y(\u_div/CryTmp[1][7] ),
	.C(FE_RN_645_0),
	.B(FE_RN_639_0),
	.A(FE_RN_629_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_750_0 (
	.Y(n57),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_749_0 (
	.Y(FE_RN_603_0),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_748_0 (
	.Y(FE_RN_602_0),
	.A(\u_div/SumTmp[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_747_0 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(FE_RN_602_0),
	.A(FE_RN_603_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_746_0 (
	.Y(FE_RN_601_0),
	.B(\u_div/BInv [4]),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_745_0 (
	.Y(FE_RN_600_0),
	.B(FE_RN_592_0),
	.A(FE_RN_601_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_744_0 (
	.Y(FE_RN_599_0),
	.C(FE_RN_574_0),
	.B(FE_RN_570_0),
	.A(FE_RN_588_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_743_0 (
	.Y(FE_RN_598_0),
	.B(FE_RN_600_0),
	.A(FE_RN_599_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_742_0 (
	.Y(\u_div/SumTmp[1][4] ),
	.B0(FE_RN_598_0),
	.A1(FE_RN_600_0),
	.A0(FE_RN_599_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_741_0 (
	.Y(FE_RN_597_0),
	.A(\u_div/BInv [4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_740_0 (
	.Y(FE_RN_596_0),
	.B(FE_RN_574_0),
	.A(FE_RN_597_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_739_0 (
	.Y(FE_RN_595_0),
	.A(FE_RN_574_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_736_0 (
	.Y(FE_RN_592_0),
	.B(FE_RN_597_0),
	.AN(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_735_0 (
	.Y(FE_RN_591_0),
	.B(quotient[2]),
	.A(\u_div/SumTmp[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M FE_RC_734_0 (
	.Y(FE_RN_590_0),
	.C0(FE_RN_573_0),
	.B0(FE_RN_591_0),
	.A1N(n37),
	.A0(quotient[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_733_0 (
	.Y(FE_RN_589_0),
	.B(FE_RN_562_0),
	.A(FE_RN_590_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_732_0 (
	.Y(FE_RN_588_0),
	.B(\u_div/CryTmp[1][2] ),
	.AN(FE_RN_589_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_731_0 (
	.Y(FE_RN_587_0),
	.B(FE_RN_570_0),
	.A(FE_RN_588_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_730_0 (
	.Y(FE_RN_586_0),
	.B(FE_RN_592_0),
	.A(FE_RN_587_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M FE_RC_728_0 (
	.Y(quotient[2]),
	.A(FE_RN_565_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_727_0 (
	.Y(FE_RN_585_0),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_726_0 (
	.Y(FE_RN_584_0),
	.B(FE_RN_585_0),
	.A(FE_RN_565_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_725_0 (
	.Y(n58),
	.B0(FE_RN_584_0),
	.A1(\u_div/SumTmp[2][1] ),
	.A0(FE_RN_565_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M FE_RC_724_0 (
	.Y(FE_RN_583_0),
	.B0(FE_RN_562_0),
	.A1N(FE_RN_572_0),
	.A0(\u_div/CryTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_723_0 (
	.Y(FE_RN_582_0),
	.A(FE_RN_562_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_722_0 (
	.Y(FE_RN_581_0),
	.A(FE_RN_572_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M FE_RC_721_0 (
	.Y(FE_RN_580_0),
	.B0(FE_RN_581_0),
	.A1N(FE_RN_582_0),
	.A0(\u_div/CryTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_720_0 (
	.Y(FE_RN_579_0),
	.B(\u_div/BInv [3]),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_719_0 (
	.Y(\u_div/SumTmp[1][3] ),
	.B1(FE_RN_579_0),
	.B0(FE_RN_580_0),
	.A1N(FE_RN_583_0),
	.A0N(FE_RN_579_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_718_0 (
	.Y(FE_RN_578_0),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(FE_RN_564_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_716_0 (
	.Y(FE_RN_576_0),
	.B(FE_RN_581_0),
	.AN(FE_RN_562_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_715_0 (
	.Y(\u_div/SumTmp[1][2] ),
	.S0(\u_div/CryTmp[1][2] ),
	.B(FE_RN_576_0),
	.A(FE_RN_578_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_714_0 (
	.Y(FE_RN_575_0),
	.A(FE_RN_572_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_713_0 (
	.Y(FE_RN_574_0),
	.B(\u_div/BInv [3]),
	.A(FE_RN_575_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_712_0 (
	.Y(FE_RN_573_0),
	.A(\u_div/BInv [3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_711_0 (
	.Y(FE_RN_572_0),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(FE_RN_564_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_710_0 (
	.Y(FE_RN_571_0),
	.B(FE_RN_573_0),
	.A(FE_RN_572_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_709_0 (
	.Y(FE_RN_570_0),
	.B(\u_div/PartRem[2][3] ),
	.A(FE_RN_571_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_707_0 (
	.Y(FE_RN_568_0),
	.A(\u_div/SumTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_705_0 (
	.Y(FE_RN_566_0),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_704_0 (
	.Y(FE_RN_565_0),
	.B(FE_RN_566_0),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_703_0 (
	.Y(FE_RN_564_0),
	.S0(FE_RN_565_0),
	.B(FE_RN_585_0),
	.A(FE_RN_568_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_702_0 (
	.Y(FE_RN_563_0),
	.A(FE_OFN11_u_div_BInv_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_701_0 (
	.Y(FE_RN_562_0),
	.B(FE_RN_563_0),
	.AN(FE_RN_564_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_675_0 (
	.Y(FE_RN_541_0),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_674_0 (
	.Y(FE_RN_540_0),
	.A(\u_div/SumTmp[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_673_0 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(n24),
	.B(FE_RN_540_0),
	.A(FE_RN_541_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_654_0 (
	.Y(FE_RN_528_0),
	.B0(FE_RN_499_0),
	.A1(FE_RN_493_0),
	.A0(FE_RN_502_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_653_0 (
	.Y(FE_RN_527_0),
	.B(\u_div/BInv [5]),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_652_0 (
	.Y(FE_RN_526_0),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_651_0 (
	.Y(FE_RN_525_0),
	.B(FE_RN_526_0),
	.AN(FE_RN_503_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_649_0 (
	.Y(FE_RN_523_0),
	.B(FE_RN_597_0),
	.AN(FE_RN_503_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_648_0 (
	.Y(FE_RN_522_0),
	.A(\u_div/CryTmp[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_647_0 (
	.Y(FE_RN_521_0),
	.C(FE_RN_522_0),
	.B(FE_RN_495_0),
	.A(FE_RN_497_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M FE_RC_646_0 (
	.Y(FE_RN_520_0),
	.D(FE_RN_493_0),
	.C(FE_RN_525_0),
	.B(FE_RN_523_0),
	.A(FE_RN_521_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_645_0 (
	.Y(FE_RN_519_0),
	.B(FE_RN_527_0),
	.A(FE_RN_520_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M FE_RC_644_0 (
	.Y(\u_div/SumTmp[2][5] ),
	.B0(FE_RN_519_0),
	.A1(FE_RN_527_0),
	.A0(FE_RN_528_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_643_0 (
	.Y(FE_RN_518_0),
	.B(\u_div/BInv [4]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_641_0 (
	.Y(FE_RN_516_0),
	.B(FE_RN_522_0),
	.A(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_640_0 (
	.Y(FE_RN_515_0),
	.B(FE_RN_503_0),
	.A(FE_RN_516_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_639_0 (
	.Y(FE_RN_514_0),
	.B(FE_RN_518_0),
	.A(FE_RN_515_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_638_0 (
	.Y(FE_RN_513_0),
	.A(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_637_0 (
	.Y(FE_RN_512_0),
	.B(FE_RN_493_0),
	.A(FE_RN_497_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_636_0 (
	.Y(FE_RN_511_0),
	.B0(FE_RN_512_0),
	.A1(FE_RN_513_0),
	.A0(FE_RN_502_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_635_0 (
	.Y(\u_div/SumTmp[2][4] ),
	.B(FE_RN_514_0),
	.A(FE_RN_511_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_633_0 (
	.Y(FE_RN_509_0),
	.B(\u_div/BInv [3]),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_632_0 (
	.Y(FE_RN_508_0),
	.B(FE_RN_522_0),
	.A(FE_RN_509_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_631_0 (
	.Y(FE_RN_507_0),
	.B(FE_RN_503_0),
	.A(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_630_0 (
	.Y(FE_RN_506_0),
	.B(\u_div/CryTmp[2][3] ),
	.A(FE_RN_507_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_629_0 (
	.Y(\u_div/SumTmp[2][3] ),
	.B(FE_RN_508_0),
	.A(FE_RN_506_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_628_0 (
	.Y(FE_RN_505_0),
	.B(\u_div/BInv [5]),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_626_0 (
	.Y(FE_RN_503_0),
	.B(FE_RN_573_0),
	.AN(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_625_0 (
	.Y(FE_RN_502_0),
	.B(\u_div/CryTmp[2][3] ),
	.A(FE_RN_503_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_624_0 (
	.Y(FE_RN_501_0),
	.C(FE_RN_502_0),
	.B(FE_RN_493_0),
	.AN(FE_RN_505_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_623_0 (
	.Y(FE_RN_500_0),
	.B(FE_RN_493_0),
	.AN(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_622_0 (
	.Y(FE_RN_499_0),
	.B(FE_RN_497_0),
	.A(FE_RN_500_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_621_0 (
	.Y(FE_RN_498_0),
	.B(\u_div/BInv [5]),
	.A(FE_RN_499_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_620_0 (
	.Y(FE_RN_497_0),
	.B(\u_div/BInv [4]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_618_0 (
	.Y(FE_RN_495_0),
	.B(\u_div/BInv [3]),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_616_0 (
	.Y(FE_RN_493_0),
	.B(FE_RN_597_0),
	.AN(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_615_0 (
	.Y(FE_RN_492_0),
	.B(FE_RN_493_0),
	.AN(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_614_0 (
	.Y(FE_RN_491_0),
	.C(FE_RN_497_0),
	.B(FE_RN_636_0),
	.A(FE_RN_492_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_613_0 (
	.Y(FE_RN_490_0),
	.B(n31),
	.A(FE_RN_491_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_612_0 (
	.Y(\u_div/CryTmp[2][6] ),
	.C(FE_RN_501_0),
	.B(FE_RN_498_0),
	.A(FE_RN_490_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_208_0 (
	.Y(n21),
	.B(n19),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_207_0 (
	.Y(FE_RN_147_0),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(FE_RN_143_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_206_0 (
	.Y(FE_RN_146_0),
	.B0(FE_RN_144_0),
	.A1N(FE_RN_143_0),
	.A0N(FE_OFN11_u_div_BInv_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_205_0 (
	.Y(FE_RN_145_0),
	.B(\u_div/CryTmp[4][2] ),
	.A(FE_RN_146_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_204_0 (
	.Y(\u_div/SumTmp[4][2] ),
	.B0(FE_RN_145_0),
	.A1(\u_div/CryTmp[4][2] ),
	.A0(FE_RN_147_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M FE_RC_203_0 (
	.Y(FE_RN_144_0),
	.C(n20),
	.B(n19),
	.AN(FE_OFN11_u_div_BInv_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_202_0 (
	.Y(FE_RN_143_0),
	.B(n20),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X8M FE_RC_201_0 (
	.Y(\u_div/CryTmp[4][3] ),
	.B1(FE_RN_143_0),
	.B0(FE_OFN11_u_div_BInv_2_),
	.A1(\u_div/CryTmp[4][2] ),
	.A0(FE_RN_144_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_97_0 (
	.Y(\u_div/PartRem[6][1] ),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_96_0 (
	.Y(FE_RN_59_0),
	.B(\u_div/CryTmp[5][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_95_0 (
	.Y(FE_RN_58_0),
	.B(FE_RN_55_0),
	.A(FE_RN_59_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_94_0 (
	.Y(\u_div/SumTmp[5][1] ),
	.B(FE_RN_58_0),
	.A(FE_RN_54_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_92_0 (
	.Y(FE_RN_56_0),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_91_0 (
	.Y(FE_RN_55_0),
	.B(FE_RN_56_0),
	.AN(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_90_0 (
	.Y(FE_RN_54_0),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_89_0 (
	.Y(FE_RN_53_0),
	.B(FE_RN_55_0),
	.A(FE_RN_54_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_88_0 (
	.Y(\u_div/CryTmp[5][2] ),
	.B(FE_RN_59_0),
	.A(FE_RN_53_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M FE_RC_77_0 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(a[6]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_76_0 (
	.Y(FE_RN_31_0),
	.B(\u_div/BInv [1]),
	.A(FE_RN_47_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_75_0 (
	.Y(\u_div/SumTmp[6][0] ),
	.B0(FE_RN_47_0),
	.A1N(a[6]),
	.A0N(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M FE_RC_74_0 (
	.Y(FE_RN_47_0),
	.B(\u_div/BInv [0]),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_72_0 (
	.Y(FE_RN_45_0),
	.B(FE_RN_31_0),
	.A(FE_RN_32_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X4M FE_RC_71_0 (
	.Y(quotient[6]),
	.C(n2),
	.B(FE_RN_33_0),
	.A(FE_RN_45_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_70_0 (
	.Y(FE_RN_44_0),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_69_0 (
	.Y(FE_RN_43_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_67_0 (
	.Y(FE_RN_41_0),
	.S0(FE_RN_56_0),
	.B(FE_RN_43_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_66_0 (
	.Y(FE_RN_40_0),
	.B(FE_RN_44_0),
	.A(FE_RN_41_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_63_0 (
	.Y(FE_RN_37_0),
	.B0(FE_RN_31_0),
	.A1N(FE_RN_56_0),
	.A0N(FE_RN_43_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_62_0 (
	.Y(FE_RN_36_0),
	.B(n1),
	.A(FE_RN_37_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_61_0 (
	.Y(\u_div/SumTmp[6][1] ),
	.B(FE_RN_40_0),
	.A(FE_RN_36_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_58_0 (
	.Y(FE_RN_33_0),
	.B(FE_RN_43_0),
	.A(FE_RN_56_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_57_0 (
	.Y(FE_RN_32_0),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X3M FE_RC_1_0 (
	.Y(\u_div/PartRem[4][2] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC11_u_div_BInv_2_ (
	.Y(FE_OFN11_u_div_BInv_2_),
	.A(\u_div/BInv [2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(\u_div/BInv [6]),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(\u_div/BInv [7]),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_3_3  (
	.S(\u_div/SumTmp[3][3] ),
	.CO(\u_div/CryTmp[3][4] ),
	.CI(\u_div/CryTmp[3][3] ),
	.B(\u_div/BInv [3]),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(\u_div/BInv [4]),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(\u_div/BInv [3]),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/PartRem[1][1] ),
	.B(\u_div/BInv [1]),
	.A(\u_div/CryTmp[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/CryTmp[1][1] ),
	.B(\u_div/PartRem[2][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(\u_div/BInv [5]),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_3_4  (
	.S(\u_div/SumTmp[3][4] ),
	.CO(\u_div/CryTmp[3][5] ),
	.CI(\u_div/CryTmp[3][4] ),
	.B(\u_div/BInv [4]),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX8M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(\u_div/PartRem[5][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX4M \u_div/u_fa_PartRem_0_5_2  (
	.S(\u_div/SumTmp[5][2] ),
	.CO(\u_div/CryTmp[5][3] ),
	.CI(\u_div/CryTmp[5][2] ),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U1 (
	.Y(n26),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U2 (
	.Y(n51),
	.B(n52),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X8M U3 (
	.Y(n67),
	.B(\u_div/BInv [3]),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U4 (
	.Y(n89),
	.B(n90),
	.A(\u_div/CryTmp[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U5 (
	.Y(n4),
	.B(\u_div/BInv [1]),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U6 (
	.Y(n68),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(quotient[5]),
	.B(n85),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U8 (
	.Y(n34),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U9 (
	.Y(n88),
	.B(b[4]),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M U10 (
	.Y(n52),
	.B(n3),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M U11 (
	.Y(\u_div/BInv [1]),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M U12 (
	.Y(n66),
	.B(n67),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U15 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(n75),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M U16 (
	.Y(n24),
	.B(n83),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U18 (
	.Y(n83),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X3M U19 (
	.Y(n1),
	.S0(n51),
	.B(\u_div/SumTmp[7][0] ),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M U20 (
	.Y(n72),
	.B(n74),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M U21 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(n66),
	.B(n65),
	.A(n196), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U23 (
	.Y(n45),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U24 (
	.Y(n5),
	.B(\u_div/CryTmp[2][1] ),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n80),
	.A(\u_div/SumTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U27 (
	.Y(n35),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U28 (
	.Y(\u_div/BInv [0]),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX6M U29 (
	.Y(\u_div/BInv [3]),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n90),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U31 (
	.Y(\u_div/BInv [2]),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(n45),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n49),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n16),
	.B(n15),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U36 (
	.Y(n18),
	.A(quotient[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M U37 (
	.Y(n87),
	.A(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(\u_div/CryTmp[4][4] ),
	.C(n12),
	.B(n13),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(n20),
	.B(quotient[5]),
	.A(\u_div/SumTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M U40 (
	.Y(\u_div/CryTmp[2][3] ),
	.C(n10),
	.B(n8),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U41 (
	.Y(n53),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U42 (
	.Y(n77),
	.B(n78),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U44 (
	.Y(n2),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U45 (
	.Y(n3),
	.B(n49),
	.A(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M U46 (
	.Y(n73),
	.B(n26),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X12M U47 (
	.Y(n82),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U48 (
	.Y(n14),
	.B(\u_div/BInv [3]),
	.A(\u_div/CryTmp[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U49 (
	.Y(n11),
	.B(\u_div/CryTmp[4][3] ),
	.A(\u_div/BInv [3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U51 (
	.Y(n9),
	.B(\u_div/CryTmp[2][2] ),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U52 (
	.Y(n10),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(\u_div/CryTmp[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U53 (
	.Y(n38),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U54 (
	.Y(n31),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M U55 (
	.Y(\u_div/CryTmp[2][2] ),
	.C(n6),
	.B(n5),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U56 (
	.Y(\u_div/SumTmp[2][1] ),
	.C(\u_div/CryTmp[2][1] ),
	.B(\u_div/BInv [1]),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2XLM U57 (
	.Y(n6),
	.B(\u_div/CryTmp[2][1] ),
	.A(\u_div/BInv [1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U58 (
	.Y(n7),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U59 (
	.Y(\u_div/SumTmp[2][2] ),
	.B(\u_div/CryTmp[2][2] ),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U60 (
	.Y(n8),
	.B(FE_OFN11_u_div_BInv_2_),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U61 (
	.Y(\u_div/SumTmp[4][3] ),
	.B(n39),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M U62 (
	.Y(n12),
	.B(\u_div/CryTmp[4][3] ),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U63 (
	.Y(n13),
	.B(\u_div/BInv [3]),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U64 (
	.Y(n48),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][1] ),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U65 (
	.Y(n85),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U66 (
	.Y(n15),
	.A(quotient[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U67 (
	.Y(n39),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U68 (
	.Y(n17),
	.B(quotient[6]),
	.A(\u_div/SumTmp[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U69 (
	.Y(n55),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U70 (
	.Y(n54),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U73 (
	.Y(n74),
	.A(\u_div/CryTmp[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U74 (
	.Y(\u_div/BInv [4]),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U75 (
	.Y(n79),
	.A(\u_div/CryTmp[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U76 (
	.Y(n76),
	.S0(n77),
	.B(\u_div/SumTmp[3][0] ),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U78 (
	.Y(n19),
	.B(n18),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(\u_div/PartRem[2][6] ),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n28),
	.A(\u_div/SumTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M U81 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(n72),
	.B(n71),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U82 (
	.Y(n81),
	.B(n83),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U84 (
	.Y(quotient[4]),
	.B(n73),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U85 (
	.Y(n37),
	.S0(n89),
	.B(n29),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U86 (
	.Y(n29),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2XLM U87 (
	.Y(n36),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U88 (
	.Y(n59),
	.S0(n81),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M U89 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(n80),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U91 (
	.Y(quotient[1]),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U94 (
	.Y(quotient[3]),
	.A(n89), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U95 (
	.Y(\u_div/PartRem[2][5] ),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U96 (
	.Y(n60),
	.A(\u_div/SumTmp[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U97 (
	.Y(n78),
	.B(\u_div/BInv [5]),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U98 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(n69),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U99 (
	.Y(n69),
	.A(\u_div/SumTmp[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U100 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(n61),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U101 (
	.Y(n61),
	.A(\u_div/SumTmp[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U103 (
	.Y(n56),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(\u_div/PartRem[2][4] ),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U105 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(n62),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n62),
	.A(\u_div/SumTmp[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U107 (
	.Y(\u_div/BInv [5]),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n70),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n71),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U111 (
	.Y(n65),
	.A(\u_div/SumTmp[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2XLM U112 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2XLM U113 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2XLM U114 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U115 (
	.Y(n75),
	.A(\u_div/SumTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U116 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n41),
	.AN(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U117 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n199),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U118 (
	.Y(n43),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U119 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(a[3]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2XLM U120 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(n60),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U121 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n42),
	.AN(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U123 (
	.Y(n42),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2XLM U124 (
	.Y(n40),
	.B(a[1]),
	.A(\u_div/BInv [0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U125 (
	.Y(n41),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U128 (
	.Y(quotient[7]),
	.B(n67),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U129 (
	.Y(\u_div/BInv [6]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U130 (
	.Y(\u_div/BInv [7]),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M U131 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(n84),
	.B(n40),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U132 (
	.Y(n91),
	.B(\u_div/CryTmp[1][7] ),
	.AN(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX4M U133 (
	.Y(n84),
	.B(b[7]),
	.AN(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_0  (
	.S(\u_div/SumTmp[4][0] ),
	.CO(\u_div/CryTmp[4][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_0  (
	.S(\u_div/SumTmp[5][0] ),
	.CO(\u_div/CryTmp[5][1] ),
	.CI(HTIE_LTIEHI_NET),
	.B(\u_div/BInv [0]),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_test_1 (
	RST, 
	TX_CLK, 
	RX_CLK, 
	RX_IN_S, 
	RX_OUT_P, 
	RX_OUT_V, 
	TX_IN_P, 
	TX_IN_V, 
	TX_OUT_S, 
	TX_OUT_V, 
	Prescale, 
	parity_enable, 
	parity_type, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_SYNC_UART_RST_M, 
	VDD, 
	VSS);
   input RST;
   input TX_CLK;
   input RX_CLK;
   input RX_IN_S;
   output [7:0] RX_OUT_P;
   output RX_OUT_V;
   input [7:0] TX_IN_P;
   input TX_IN_V;
   output TX_OUT_S;
   output TX_OUT_V;
   input [5:0] Prescale;
   input parity_enable;
   input parity_type;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_SYNC_UART_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n4;

   // Module instantiations
   UART_TX_test_1 U0_UART_TX (
	.P_DATA({ TX_IN_P[7],
		TX_IN_P[6],
		TX_IN_P[5],
		TX_IN_P[4],
		TX_IN_P[3],
		TX_IN_P[2],
		TX_IN_P[1],
		TX_IN_P[0] }),
	.Data_Valid(TX_IN_V),
	.PAR_EN(parity_enable),
	.PAR_TYP(parity_type),
	.CLK(TX_CLK),
	.RST(RST),
	.TX_OUT(TX_OUT_S),
	.busy(TX_OUT_V),
	.test_si(n4),
	.test_so(test_so),
	.test_se(test_se),
	.FE_OFN3_SYNC_UART_RST_M(FE_OFN3_SYNC_UART_RST_M), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_RX_test_1 U0_UART_RX (
	.RX_IN(RX_IN_S),
	.PAR_EN(parity_enable),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.PAR_TYP(parity_type),
	.RX_CLK(RX_CLK),
	.RST(FE_OFN3_SYNC_UART_RST_M),
	.P_DATA({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.data_Valid(RX_OUT_V),
	.test_si(test_si),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TX_test_1 (
	P_DATA, 
	Data_Valid, 
	PAR_EN, 
	PAR_TYP, 
	CLK, 
	RST, 
	TX_OUT, 
	busy, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_SYNC_UART_RST_M, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input Data_Valid;
   input PAR_EN;
   input PAR_TYP;
   input CLK;
   input RST;
   output TX_OUT;
   output busy;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_SYNC_UART_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire ser_done;
   wire ser_en;
   wire par_bit;
   wire ser_data;
   wire n4;
   wire [1:0] mux_sel;

   // Module instantiations
   tx_controller_test_1 U1 (
	.Data_Valid(Data_Valid),
	.PAR_EN(PAR_EN),
	.ser_done(ser_done),
	.CLK(CLK),
	.RST(FE_OFN3_SYNC_UART_RST_M),
	.ser_en(ser_en),
	.mux_sel({ mux_sel[1],
		mux_sel[0] }),
	.busy(busy),
	.test_si(n4),
	.test_so(test_so),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   Parity_Calc_test_1 P1 (
	.CLK(CLK),
	.RST(RST),
	.PAR_EN(PAR_EN),
	.PAR_TYP(PAR_TYP),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.busy(busy),
	.Data_Valid(Data_Valid),
	.par_bit(par_bit),
	.test_si(test_si),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   Serializer_test_1 S1 (
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.Data_Valid(Data_Valid),
	.busy(busy),
	.ser_en(ser_en),
	.CLK(CLK),
	.RST(RST),
	.ser_data(ser_data),
	.ser_done(ser_done),
	.test_si(par_bit),
	.test_so(n4),
	.test_se(test_se),
	.FE_OFN3_SYNC_UART_RST_M(FE_OFN3_SYNC_UART_RST_M), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_4_1 M1 (
	.A(1'b0),
	.B(ser_data),
	.C(par_bit),
	.D(1'b1),
	.sel({ mux_sel[1],
		mux_sel[0] }),
	.out(TX_OUT), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module tx_controller_test_1 (
	Data_Valid, 
	PAR_EN, 
	ser_done, 
	CLK, 
	RST, 
	ser_en, 
	mux_sel, 
	busy, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input Data_Valid;
   input PAR_EN;
   input ser_done;
   input CLK;
   input RST;
   output ser_en;
   output [1:0] mux_sel;
   output busy;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n5),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n6),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U6 (
	.Y(mux_sel[1]),
	.B0(n12),
	.A1(n5),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n12),
	.B(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI33X2M U8 (
	.Y(ser_en),
	.B2(current_state[0]),
	.B1(ser_done),
	.B0(n10),
	.A2(current_state[1]),
	.A1(current_state[2]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n10),
	.B(n7),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n5),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n7),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U12 (
	.Y(busy),
	.C0(n10),
	.B1(n5),
	.B0(current_state[2]),
	.A1(n7),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U13 (
	.Y(next_state[1]),
	.B0(n4),
	.A2(n10),
	.A1(current_state[0]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n4),
	.A(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(next_state[0]),
	.C(current_state[0]),
	.B(current_state[2]),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U16 (
	.Y(n11),
	.B1(n6),
	.B0(Data_Valid),
	.A2(PAR_EN),
	.A1(current_state[1]),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(next_state[2]),
	.B(n10),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U18 (
	.Y(n9),
	.B0(current_state[0]),
	.A1(n8),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n6),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n8),
	.A(PAR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U21 (
	.Y(mux_sel[0]),
	.B0(n12),
	.A1(current_state[0]),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Parity_Calc_test_1 (
	CLK, 
	RST, 
	PAR_EN, 
	PAR_TYP, 
	P_DATA, 
	busy, 
	Data_Valid, 
	par_bit, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input PAR_EN;
   input PAR_TYP;
   input [7:0] P_DATA;
   input busy;
   input Data_Valid;
   output par_bit;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;

   // Module instantiations
   SDFFRQX2M par_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(par_bit),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(n5),
	.B(P_DATA[2]),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U3 (
	.Y(n3),
	.C(n6),
	.B(P_DATA[4]),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(n6),
	.B(P_DATA[6]),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U5 (
	.Y(n8),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(par_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U6 (
	.Y(n2),
	.C(PAR_EN),
	.B(Data_Valid),
	.AN(busy), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U7 (
	.Y(n1),
	.C(n4),
	.B(PAR_TYP),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n4),
	.C(n5),
	.B(P_DATA[0]),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Serializer_test_1 (
	P_DATA, 
	Data_Valid, 
	busy, 
	ser_en, 
	CLK, 
	RST, 
	ser_data, 
	ser_done, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN3_SYNC_UART_RST_M, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input Data_Valid;
   input busy;
   input ser_en;
   input CLK;
   input RST;
   output ser_data;
   output ser_done;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN3_SYNC_UART_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n17;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n15;
   wire n16;
   wire n18;
   wire n48;
   wire n49;
   wire n52;
   wire n53;
   wire [7:0] temp_data;
   wire [3:0] count;

   assign test_so = temp_data[7] ;

   // Module instantiations
   SDFFRQX2M \temp_data_reg[6]  (
	.SI(temp_data[5]),
	.SE(n53),
	.RN(FE_OFN3_SYNC_UART_RST_M),
	.Q(temp_data[6]),
	.D(n38),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[5]  (
	.SI(temp_data[4]),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[5]),
	.D(n39),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[4]  (
	.SI(temp_data[3]),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[4]),
	.D(n40),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[3]  (
	.SI(temp_data[2]),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[3]),
	.D(n41),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[2]  (
	.SI(temp_data[1]),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[2]),
	.D(n42),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[1]  (
	.SI(temp_data[0]),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[1]),
	.D(n43),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[0]  (
	.SI(ser_data),
	.SE(n53),
	.RN(RST),
	.Q(temp_data[0]),
	.D(n44),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M ser_data_reg (
	.SI(n49),
	.SE(n53),
	.RN(RST),
	.Q(ser_data),
	.D(n36),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \temp_data_reg[7]  (
	.SI(temp_data[6]),
	.SE(n53),
	.RN(FE_OFN3_SYNC_UART_RST_M),
	.Q(temp_data[7]),
	.D(n37),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[2]  (
	.SI(count[1]),
	.SE(n53),
	.RN(RST),
	.Q(count[2]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[0]  (
	.SI(test_si),
	.SE(n53),
	.RN(RST),
	.Q(count[0]),
	.D(n47),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \count_reg[1]  (
	.SI(count[0]),
	.SE(n53),
	.RN(RST),
	.Q(count[1]),
	.D(n45),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \count_reg[3]  (
	.SI(n48),
	.SE(n53),
	.RN(RST),
	.QN(n17),
	.Q(n49),
	.D(n46),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U17 (
	.Y(ser_done),
	.D(count[2]),
	.C(count[1]),
	.B(count[0]),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(n19),
	.B(n21),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(n20),
	.B(n19),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n16),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U21 (
	.Y(n35),
	.B(ser_done),
	.AN(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n18),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U23 (
	.Y(n21),
	.B(busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U24 (
	.Y(n31),
	.B1(ser_en),
	.B0(n16),
	.A1N(n16),
	.A0N(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U25 (
	.Y(n45),
	.B1(n32),
	.B0(count[1]),
	.A1N(count[1]),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U26 (
	.Y(n30),
	.B0(n31),
	.A1(n16),
	.A0(count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U27 (
	.Y(n46),
	.B0(n34),
	.A1(n17),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U28 (
	.Y(n34),
	.D(n17),
	.C(n18),
	.B(count[1]),
	.A(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U29 (
	.Y(n33),
	.B0(n30),
	.A1(n48),
	.A0(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U30 (
	.Y(n32),
	.B(n35),
	.A(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(n47),
	.B(n16),
	.A(count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n15),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U33 (
	.Y(n29),
	.B1(count[2]),
	.B0(n30),
	.A2(n18),
	.A1(n48),
	.A0(count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U34 (
	.Y(n44),
	.B0(n28),
	.A1N(n20),
	.A0N(temp_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U35 (
	.Y(n28),
	.B1(n21),
	.B0(P_DATA[0]),
	.A1(n19),
	.A0(temp_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U36 (
	.Y(n43),
	.B0(n27),
	.A1N(temp_data[1]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U37 (
	.Y(n27),
	.B1(n21),
	.B0(P_DATA[1]),
	.A1(n19),
	.A0(temp_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U38 (
	.Y(n42),
	.B0(n26),
	.A1N(temp_data[2]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U39 (
	.Y(n26),
	.B1(n21),
	.B0(P_DATA[2]),
	.A1(n19),
	.A0(temp_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U40 (
	.Y(n41),
	.B0(n25),
	.A1N(temp_data[3]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U41 (
	.Y(n25),
	.B1(n21),
	.B0(P_DATA[3]),
	.A1(n19),
	.A0(temp_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U42 (
	.Y(n40),
	.B0(n24),
	.A1N(temp_data[4]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U43 (
	.Y(n24),
	.B1(n21),
	.B0(P_DATA[4]),
	.A1(n19),
	.A0(temp_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U44 (
	.Y(n39),
	.B0(n23),
	.A1N(temp_data[5]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U45 (
	.Y(n23),
	.B1(n21),
	.B0(P_DATA[5]),
	.A1(n19),
	.A0(temp_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U46 (
	.Y(n38),
	.B0(n22),
	.A1N(temp_data[6]),
	.A0N(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U47 (
	.Y(n22),
	.B1(n21),
	.B0(P_DATA[6]),
	.A1(n19),
	.A0(temp_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U48 (
	.Y(n36),
	.B1(n20),
	.B0(ser_data),
	.A1(temp_data[0]),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U49 (
	.Y(n37),
	.B1(n21),
	.B0(P_DATA[7]),
	.A1(temp_data[7]),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n48),
	.A(count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U51 (
	.Y(n52),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U52 (
	.Y(n53),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_4_1 (
	A, 
	B, 
	C, 
	D, 
	sel, 
	out, 
	VDD, 
	VSS);
   input A;
   input B;
   input C;
   input D;
   input [1:0] sel;
   output out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire n2;
   wire n3;
   wire n1;
   wire n4;
   wire n5;
   wire n6;
   wire n7;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U1 (
	.Y(out),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(n4),
	.A(sel[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U3 (
	.Y(n5),
	.B(n3),
	.A(sel[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U4 (
	.Y(n6),
	.B(n4),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U5 (
	.Y(n1),
	.B(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U6 (
	.Y(n3),
	.B1(B),
	.B0(sel[0]),
	.A1(n7),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U7 (
	.Y(n2),
	.B1(sel[0]),
	.B0(HTIE_LTIEHI_NET),
	.A1(n7),
	.A0(C), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n7),
	.A(sel[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_test_1 (
	RX_IN, 
	PAR_EN, 
	Prescale, 
	PAR_TYP, 
	RX_CLK, 
	RST, 
	P_DATA, 
	data_Valid, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input RX_IN;
   input PAR_EN;
   input [5:0] Prescale;
   input PAR_TYP;
   input RX_CLK;
   input RST;
   output [7:0] P_DATA;
   output data_Valid;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire samp_en;
   wire sampled_bit;
   wire cnt_en;
   wire stp_err;
   wire strt_glitch;
   wire par_err;
   wire par_chk_en;
   wire strt_chk_en;
   wire stp_chk_en;
   wire deser_en;
   wire n3;
   wire n4;
   wire n5;
   wire [2:0] edge_cnt;
   wire [3:0] bit_cnt;

   assign test_so = strt_glitch ;

   // Module instantiations
   data_sampling_test_1 D0 (
	.RX_IN(RX_IN),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.enable(samp_en),
	.edge_count({ edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.CLK(RX_CLK),
	.RST(RST),
	.sampled_bit(sampled_bit),
	.test_si(test_si),
	.test_so(n5),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   edge_bit_counter_test_1 E_B_c (
	.enable(cnt_en),
	.CLK(RX_CLK),
	.RST(RST),
	.bit_cnt({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }),
	.edge_cnt({ edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.test_si(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   RX_controller_test_1 RX0 (
	.RX_IN(RX_IN),
	.PAR_EN(PAR_EN),
	.edge_cnt({ edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.bit_cnt({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }),
	.stp_err(stp_err),
	.strt_glitch(strt_glitch),
	.par_err(par_err),
	.CLK(RX_CLK),
	.RST(RST),
	.par_chk_en(par_chk_en),
	.strt_chk_en(strt_chk_en),
	.stp_chk_en(stp_chk_en),
	.deser_en(deser_en),
	.samp_en(samp_en),
	.cnt_en(cnt_en),
	.data_valid(data_Valid),
	.test_so(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   stop_check_test_1 STP0 (
	.sampled_bit(sampled_bit),
	.enable(stp_chk_en),
	.CLK(RX_CLK),
	.RST(RST),
	.stp_err(stp_err),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   strt_check_test_1 STR0 (
	.enable(strt_chk_en),
	.sampled_bit(sampled_bit),
	.CLK(RX_CLK),
	.RST(RST),
	.strt_glitch(strt_glitch),
	.test_si(stp_err),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_check_test_1 Par0 (
	.enable(par_chk_en),
	.sampled_bit(sampled_bit),
	.PAR_TYP(PAR_TYP),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.CLK(RX_CLK),
	.RST(RST),
	.par_err(par_err),
	.test_si(edge_cnt[2]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_test_1 DSR0 (
	.sampled_bit(sampled_bit),
	.edge_cnt({ edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }),
	.enable(deser_en),
	.CLK(RX_CLK),
	.RST(RST),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.test_si(n5),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_test_1 (
	RX_IN, 
	Prescale, 
	enable, 
	edge_count, 
	CLK, 
	RST, 
	sampled_bit, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input RX_IN;
   input [5:0] Prescale;
   input enable;
   input [2:0] edge_count;
   input CLK;
   input RST;
   output sampled_bit;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \half_minus_one[0] ;
   wire n12;
   wire n13;
   wire n14;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n8;

   assign \half_minus_one[0]  = Prescale[1] ;

   // Module instantiations
   SDFFRX1M \sample_test_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.QN(n14),
	.Q(n8),
	.D(n30),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \sample_test_reg[1]  (
	.SI(n8),
	.SE(test_se),
	.RN(RST),
	.QN(n13),
	.Q(n7),
	.D(n31),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \sample_test_reg[2]  (
	.SI(n7),
	.SE(test_se),
	.RN(RST),
	.QN(n12),
	.Q(test_so),
	.D(n32),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U7 (
	.Y(sampled_bit),
	.B0(n13),
	.A1(n12),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U8 (
	.Y(n30),
	.B1(n20),
	.B0(n19),
	.A2(n2),
	.A1(n3),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n2),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n3),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U11 (
	.Y(n20),
	.C(n23),
	.B(n22),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U12 (
	.Y(n31),
	.B1(n25),
	.B0(n13),
	.A1N(n25),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U13 (
	.Y(n25),
	.B0(enable),
	.A2(n26),
	.A1(n4),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n4),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U15 (
	.Y(n26),
	.C(n5),
	.B(Prescale[3]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U16 (
	.Y(n32),
	.B1(n12),
	.B0(n28),
	.A1N(n28),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U17 (
	.Y(n28),
	.B0(enable),
	.A2(n27),
	.A1(n21),
	.A0(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(n29),
	.B(Prescale[3]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U19 (
	.Y(n23),
	.C(n24),
	.B(Prescale[3]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U20 (
	.Y(n24),
	.B(n5),
	.AN(\half_minus_one[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U21 (
	.Y(n22),
	.C(Prescale[2]),
	.B(edge_count[1]),
	.A(\half_minus_one[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(n19),
	.B(enable),
	.A(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n21),
	.B(edge_count[0]),
	.A(\half_minus_one[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U24 (
	.Y(n27),
	.B(Prescale[2]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n5),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_test_1 (
	enable, 
	CLK, 
	RST, 
	bit_cnt, 
	edge_cnt, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input enable;
   input CLK;
   input RST;
   output [3:0] bit_cnt;
   output [2:0] edge_cnt;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n8;
   wire n9;
   wire n10;
   wire n11;

   // Module instantiations
   SDFFRQX2M \bit_cnt_reg[3]  (
	.SI(bit_cnt[2]),
	.SE(test_se),
	.RN(RST),
	.Q(bit_cnt[3]),
	.D(n28),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_reg[2]  (
	.SI(n9),
	.SE(test_se),
	.RN(RST),
	.Q(bit_cnt[2]),
	.D(n23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_reg[2]  (
	.SI(n8),
	.SE(test_se),
	.RN(RST),
	.Q(edge_cnt[2]),
	.D(n27),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_reg[0]  (
	.SI(n11),
	.SE(test_se),
	.RN(RST),
	.Q(edge_cnt[0]),
	.D(n26),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_reg[1]  (
	.SI(edge_cnt[0]),
	.SE(test_se),
	.RN(RST),
	.Q(edge_cnt[1]),
	.D(n25),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(bit_cnt[0]),
	.D(n29),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_reg[1]  (
	.SI(bit_cnt[0]),
	.SE(test_se),
	.RN(RST),
	.Q(bit_cnt[1]),
	.D(n24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U10 (
	.Y(n17),
	.B0(enable),
	.A1(n20),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U11 (
	.Y(n22),
	.B(n19),
	.AN(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U12 (
	.Y(n13),
	.B(n9),
	.AN(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U13 (
	.Y(n28),
	.B1(n11),
	.B0(n13),
	.A2(n10),
	.A1(n12),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n21),
	.B(n11),
	.A(bit_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n11),
	.A(bit_cnt[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U16 (
	.Y(n23),
	.B1(n10),
	.B0(n13),
	.A2(n9),
	.A1(bit_cnt[2]),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U17 (
	.Y(n25),
	.B1(n16),
	.B0(edge_cnt[1]),
	.A1(n8),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U18 (
	.Y(n24),
	.B1(n12),
	.B0(bit_cnt[1]),
	.A1(n9),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U19 (
	.Y(n16),
	.C(n19),
	.B(edge_cnt[0]),
	.AN(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U20 (
	.Y(n26),
	.B(n17),
	.A(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U21 (
	.Y(n20),
	.D(n10),
	.C(bit_cnt[0]),
	.B(bit_cnt[1]),
	.A(bit_cnt[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U22 (
	.Y(n19),
	.C(edge_cnt[2]),
	.B(edge_cnt[0]),
	.A(edge_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U23 (
	.Y(n15),
	.B(n17),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U24 (
	.Y(n12),
	.C(n22),
	.B(n20),
	.A(bit_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U25 (
	.Y(n27),
	.B0(n18),
	.A1(n16),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U26 (
	.Y(n18),
	.B0(edge_cnt[2]),
	.A1N(n15),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n9),
	.A(bit_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n10),
	.A(bit_cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n14),
	.B(bit_cnt[0]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n29),
	.B(n22),
	.A(bit_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n8),
	.A(edge_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RX_controller_test_1 (
	RX_IN, 
	PAR_EN, 
	edge_cnt, 
	bit_cnt, 
	stp_err, 
	strt_glitch, 
	par_err, 
	CLK, 
	RST, 
	par_chk_en, 
	strt_chk_en, 
	stp_chk_en, 
	deser_en, 
	samp_en, 
	cnt_en, 
	data_valid, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input RX_IN;
   input PAR_EN;
   input [2:0] edge_cnt;
   input [3:0] bit_cnt;
   input stp_err;
   input strt_glitch;
   input par_err;
   input CLK;
   input RST;
   output par_chk_en;
   output strt_chk_en;
   output stp_chk_en;
   output deser_en;
   output samp_en;
   output cnt_en;
   output data_valid;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n10;
   wire n11;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = n8 ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[0]  (
	.SI(par_err),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[2]  (
	.SI(n7),
	.SE(test_se),
	.RN(RST),
	.QN(n8),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n22),
	.B(n6),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U8 (
	.Y(stp_chk_en),
	.B(n11),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n11),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(cnt_en),
	.B(n22),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(deser_en),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(n16),
	.B(current_state[2]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U14 (
	.Y(n19),
	.B1(par_chk_en),
	.B0(par_err),
	.A1(n10),
	.A0(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U15 (
	.Y(next_state[2]),
	.B0(n14),
	.A2(n13),
	.A1(par_err),
	.A0(par_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U16 (
	.Y(next_state[1]),
	.B0(n15),
	.A2(n13),
	.A1(strt_glitch),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U17 (
	.Y(n15),
	.B0(deser_en),
	.A2(n16),
	.A1(n5),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n5),
	.A(par_err), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U19 (
	.Y(data_valid),
	.C(n8),
	.B(current_state[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U20 (
	.Y(n13),
	.C(edge_cnt[2]),
	.B(edge_cnt[0]),
	.A(edge_cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U21 (
	.Y(n14),
	.C(n9),
	.B(stp_chk_en),
	.AN(stp_err), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n9),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U23 (
	.Y(n10),
	.C(current_state[0]),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U24 (
	.Y(samp_en),
	.B(n11),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U26 (
	.Y(par_chk_en),
	.B(current_state[0]),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n6),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U28 (
	.Y(n20),
	.B0(data_valid),
	.A1N(current_state[2]),
	.A0N(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U29 (
	.Y(next_state[0]),
	.C(n18),
	.B(n14),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U30 (
	.Y(n17),
	.D(n21),
	.C(bit_cnt[3]),
	.B(deser_en),
	.A(PAR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U31 (
	.Y(n18),
	.B1(n13),
	.B0(n19),
	.A1N(n20),
	.A0N(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U32 (
	.Y(n21),
	.D(n13),
	.C(bit_cnt[0]),
	.B(bit_cnt[1]),
	.A(bit_cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(strt_chk_en),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \current_state_reg[1]  (
	.SI(n6),
	.SE(test_se),
	.RN(RST),
	.QN(n7),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stop_check_test_1 (
	sampled_bit, 
	enable, 
	CLK, 
	RST, 
	stp_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input sampled_bit;
   input enable;
   input CLK;
   input RST;
   output stp_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire n1;

   // Module instantiations
   SDFFRQX2M stp_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(stp_err),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U2 (
	.Y(n3),
	.B1(n1),
	.B0(sampled_bit),
	.A1N(n1),
	.A0N(stp_err), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n1),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module strt_check_test_1 (
	enable, 
	sampled_bit, 
	CLK, 
	RST, 
	strt_glitch, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input enable;
   input sampled_bit;
   input CLK;
   input RST;
   output strt_glitch;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;

   // Module instantiations
   SDFFRQX2M strt_glitch_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(strt_glitch),
	.D(n2),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U2 (
	.Y(n2),
	.B1(enable),
	.B0(sampled_bit),
	.A1N(enable),
	.A0(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_check_test_1 (
	enable, 
	sampled_bit, 
	PAR_TYP, 
	P_DATA, 
	CLK, 
	RST, 
	par_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input enable;
   input sampled_bit;
   input PAR_TYP;
   input [7:0] P_DATA;
   input CLK;
   input RST;
   output par_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire par_bit;
   wire N9;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;

   // Module instantiations
   SDFFRQX2M par_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(par_bit),
	.D(N9),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M par_err_reg (
	.SI(par_bit),
	.SE(test_se),
	.RN(RST),
	.Q(par_err),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(n6),
	.B(P_DATA[6]),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U4 (
	.Y(N9),
	.C(n4),
	.B(n3),
	.A(PAR_TYP), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U5 (
	.Y(n4),
	.C(n5),
	.B(P_DATA[0]),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U6 (
	.Y(n3),
	.C(n6),
	.B(P_DATA[4]),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n5),
	.B(P_DATA[2]),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U8 (
	.Y(n8),
	.B1(enable),
	.B0(n1),
	.A1N(enable),
	.A0N(par_err), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n1),
	.B(par_bit),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_test_1 (
	sampled_bit, 
	edge_cnt, 
	enable, 
	CLK, 
	RST, 
	P_DATA, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input sampled_bit;
   input [2:0] edge_cnt;
   input enable;
   input CLK;
   input RST;
   output [7:0] P_DATA;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n4;
   wire n5;
   wire n8;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n32;
   wire n34;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n3;
   wire n6;
   wire n7;
   wire n9;
   wire [2:0] cnt;

   assign test_so = cnt[2] ;

   // Module instantiations
   SDFFRQX2M \P_DATA_reg[5]  (
	.SI(P_DATA[4]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[5]),
	.D(n39),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[1]  (
	.SI(P_DATA[0]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[1]),
	.D(n43),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[4]  (
	.SI(P_DATA[3]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[4]),
	.D(n40),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[0]),
	.D(n44),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[7]  (
	.SI(P_DATA[6]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[7]),
	.D(n37),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[3]  (
	.SI(P_DATA[2]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[3]),
	.D(n41),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[6]  (
	.SI(P_DATA[5]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[6]),
	.D(n38),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[2]  (
	.SI(P_DATA[1]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[2]),
	.D(n42),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cnt_reg[2]  (
	.SI(cnt[1]),
	.SE(test_se),
	.RN(RST),
	.Q(cnt[2]),
	.D(n32),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cnt_reg[1]  (
	.SI(n3),
	.SE(test_se),
	.RN(RST),
	.Q(cnt[1]),
	.D(n34),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cnt_reg[0]  (
	.SI(P_DATA[7]),
	.SE(test_se),
	.RN(RST),
	.Q(cnt[0]),
	.D(n36),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n17),
	.B(n22),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n9),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U5 (
	.Y(n10),
	.B(sampled_bit),
	.AN(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n7),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U7 (
	.Y(n34),
	.C0(n8),
	.B1(n6),
	.B0(n9),
	.A1(n5),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U8 (
	.Y(n36),
	.B(n9),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n15),
	.B(n3),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U10 (
	.Y(n4),
	.D(edge_cnt[2]),
	.C(enable),
	.B(edge_cnt[1]),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(n22),
	.B(cnt[2]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U12 (
	.Y(n32),
	.B1(n7),
	.B0(n2),
	.A1N(cnt[2]),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U13 (
	.Y(n1),
	.B(n4),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n12),
	.B(n9),
	.A(cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U15 (
	.Y(n41),
	.B0(n18),
	.A1(n17),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U16 (
	.Y(n18),
	.B0(P_DATA[3]),
	.A1(n7),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n37),
	.B0(n11),
	.A1(n10),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U18 (
	.Y(n11),
	.B0(P_DATA[7]),
	.A1(n12),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U19 (
	.Y(n42),
	.B0(n19),
	.A1(n17),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U20 (
	.Y(n19),
	.B0(P_DATA[2]),
	.A1(n8),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U21 (
	.Y(n44),
	.B0(n21),
	.A1(n17),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U22 (
	.Y(n21),
	.B0(P_DATA[0]),
	.A1(n15),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U23 (
	.Y(n43),
	.B0(n20),
	.A1(n17),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U24 (
	.Y(n20),
	.B0(P_DATA[1]),
	.A1(n5),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U25 (
	.Y(n39),
	.B0(n14),
	.A1(n10),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U26 (
	.Y(n14),
	.B0(P_DATA[5]),
	.A1(n12),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U27 (
	.Y(n38),
	.B0(n13),
	.A1(n8),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U28 (
	.Y(n13),
	.B0(P_DATA[6]),
	.A1(n8),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U29 (
	.Y(n40),
	.B0(n16),
	.A1(n15),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U30 (
	.Y(n16),
	.B0(P_DATA[4]),
	.A1(n15),
	.A0(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n2),
	.B(cnt[0]),
	.A(cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n8),
	.B(n3),
	.A(cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U33 (
	.Y(n5),
	.B(n6),
	.A(cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n3),
	.A(cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U35 (
	.Y(n6),
	.A(cnt[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Asynch_FIFO_test_1 (
	winc, 
	wclk, 
	wrst_n, 
	rinc, 
	rclk, 
	rrst_n, 
	wdata, 
	rdata, 
	wfull, 
	rempty, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_SYNC_REF_RST_M, 
	VDD, 
	VSS);
   input winc;
   input wclk;
   input wrst_n;
   input rinc;
   input rclk;
   input rrst_n;
   input [7:0] wdata;
   output [7:0] rdata;
   output wfull;
   output rempty;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_SYNC_REF_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire [3:0] g_rptr;
   wire [3:0] wq2_rptr;
   wire [3:0] g_wptr;
   wire [3:0] rq2_wptr;
   wire [2:0] waddr;
   wire [2:0] raddr;

   assign test_so1 = wq2_rptr[3] ;
   assign test_so2 = g_wptr[3] ;

   // Module instantiations
   BIT_SYNC_NUM_STAGES2_BUS_WIDTH4_test_0 u_r2w_sync (
	.CLK(wclk),
	.RST(wrst_n),
	.ASYNC({ g_rptr[3],
		g_rptr[2],
		g_rptr[1],
		g_rptr[0] }),
	.SYNC({ wq2_rptr[3],
		wq2_rptr[2],
		wq2_rptr[1],
		wq2_rptr[0] }),
	.test_se(test_se),
	.FE_OFN0_SYNC_REF_RST_M(FE_OFN0_SYNC_REF_RST_M), 
	.VDD(VDD), 
	.VSS(VSS));
   BIT_SYNC_NUM_STAGES2_BUS_WIDTH4_test_1 u_w2r_sync (
	.CLK(rclk),
	.RST(rrst_n),
	.ASYNC({ g_wptr[3],
		g_wptr[2],
		g_wptr[1],
		g_wptr[0] }),
	.SYNC({ rq2_wptr[3],
		rq2_wptr[2],
		rq2_wptr[1],
		rq2_wptr[0] }),
	.test_si(test_si2),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_mem_Data_Width8_DEPTH8_POI_SIZE4_test_1 fifomem (
	.wclk(wclk),
	.wrst_n(wrst_n),
	.winc(winc),
	.wfull(wfull),
	.wdata({ wdata[7],
		wdata[6],
		wdata[5],
		wdata[4],
		wdata[3],
		wdata[2],
		wdata[1],
		wdata[0] }),
	.waddr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.raddr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.rdata({ rdata[7],
		rdata[6],
		rdata[5],
		rdata[4],
		rdata[3],
		rdata[2],
		rdata[1],
		rdata[0] }),
	.test_si(test_si1),
	.test_so(n3),
	.test_se(test_se),
	.FE_OFN0_SYNC_REF_RST_M(FE_OFN0_SYNC_REF_RST_M), 
	.VDD(VDD), 
	.VSS(VSS));
   r_empty_P_SIZE4_test_1 rptr_empty (
	.rinc(rinc),
	.rclk(rclk),
	.rrst_n(rrst_n),
	.rq2_wptr({ rq2_wptr[3],
		rq2_wptr[2],
		rq2_wptr[1],
		rq2_wptr[0] }),
	.rempty(rempty),
	.raddr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.g_rptr({ g_rptr[3],
		g_rptr[2],
		g_rptr[1],
		g_rptr[0] }),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   w_full_POI_SIZE4_test_1 wptr_full (
	.winc(winc),
	.wclk(wclk),
	.wrst_n(wrst_n),
	.wq2_rptr({ wq2_rptr[3],
		wq2_rptr[2],
		wq2_rptr[1],
		wq2_rptr[0] }),
	.wfull(wfull),
	.waddr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.g_wptr({ g_wptr[3],
		g_wptr[2],
		g_wptr[1],
		g_wptr[0] }),
	.test_si(rq2_wptr[3]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module BIT_SYNC_NUM_STAGES2_BUS_WIDTH4_test_0 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_se, 
	FE_OFN0_SYNC_REF_RST_M, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [3:0] ASYNC;
   output [3:0] SYNC;
   input test_se;
   input FE_OFN0_SYNC_REF_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \sync_reg[3][0] ;
   wire \sync_reg[2][0] ;
   wire \sync_reg[1][0] ;
   wire \sync_reg[0][0] ;

   // Module instantiations
   SDFFRQX2M \sync_reg_reg[3][1]  (
	.SI(\sync_reg[3][0] ),
	.SE(test_se),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(SYNC[3]),
	.D(\sync_reg[3][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[2][1]  (
	.SI(\sync_reg[2][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[2]),
	.D(\sync_reg[2][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[1][1]  (
	.SI(\sync_reg[1][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[1]),
	.D(\sync_reg[1][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0][1]  (
	.SI(\sync_reg[0][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[0]),
	.D(\sync_reg[0][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[3][0]  (
	.SI(SYNC[2]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[3][0] ),
	.D(ASYNC[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[2][0]  (
	.SI(SYNC[1]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[2][0] ),
	.D(ASYNC[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[1][0]  (
	.SI(SYNC[0]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[1][0] ),
	.D(ASYNC[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0][0]  (
	.SI(ASYNC[3]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[0][0] ),
	.D(ASYNC[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module BIT_SYNC_NUM_STAGES2_BUS_WIDTH4_test_1 (
	CLK, 
	RST, 
	ASYNC, 
	SYNC, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [3:0] ASYNC;
   output [3:0] SYNC;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \sync_reg[3][0] ;
   wire \sync_reg[2][0] ;
   wire \sync_reg[1][0] ;
   wire \sync_reg[0][0] ;

   // Module instantiations
   SDFFRQX2M \sync_reg_reg[2][1]  (
	.SI(\sync_reg[2][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[2]),
	.D(\sync_reg[2][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[1][1]  (
	.SI(\sync_reg[1][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[1]),
	.D(\sync_reg[1][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0][1]  (
	.SI(\sync_reg[0][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[0]),
	.D(\sync_reg[0][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[3][0]  (
	.SI(SYNC[2]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[3][0] ),
	.D(ASYNC[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[2][0]  (
	.SI(SYNC[1]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[2][0] ),
	.D(ASYNC[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[1][0]  (
	.SI(SYNC[0]),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[1][0] ),
	.D(ASYNC[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0][0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\sync_reg[0][0] ),
	.D(ASYNC[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \sync_reg_reg[3][1]  (
	.SI(\sync_reg[3][0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC[3]),
	.D(\sync_reg[3][0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_mem_Data_Width8_DEPTH8_POI_SIZE4_test_1 (
	wclk, 
	wrst_n, 
	winc, 
	wfull, 
	wdata, 
	waddr, 
	raddr, 
	rdata, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN0_SYNC_REF_RST_M, 
	VDD, 
	VSS);
   input wclk;
   input wrst_n;
   input winc;
   input wfull;
   input [7:0] wdata;
   input [2:0] waddr;
   input [2:0] raddr;
   output [7:0] rdata;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN0_SYNC_REF_RST_M;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N9;
   wire N10;
   wire N11;
   wire \MEM[7][7] ;
   wire \MEM[7][6] ;
   wire \MEM[7][5] ;
   wire \MEM[7][4] ;
   wire \MEM[7][3] ;
   wire \MEM[7][2] ;
   wire \MEM[7][1] ;
   wire \MEM[7][0] ;
   wire \MEM[6][7] ;
   wire \MEM[6][6] ;
   wire \MEM[6][5] ;
   wire \MEM[6][4] ;
   wire \MEM[6][3] ;
   wire \MEM[6][2] ;
   wire \MEM[6][1] ;
   wire \MEM[6][0] ;
   wire \MEM[5][7] ;
   wire \MEM[5][6] ;
   wire \MEM[5][5] ;
   wire \MEM[5][4] ;
   wire \MEM[5][3] ;
   wire \MEM[5][2] ;
   wire \MEM[5][1] ;
   wire \MEM[5][0] ;
   wire \MEM[4][7] ;
   wire \MEM[4][6] ;
   wire \MEM[4][5] ;
   wire \MEM[4][4] ;
   wire \MEM[4][3] ;
   wire \MEM[4][2] ;
   wire \MEM[4][1] ;
   wire \MEM[4][0] ;
   wire \MEM[3][7] ;
   wire \MEM[3][6] ;
   wire \MEM[3][5] ;
   wire \MEM[3][4] ;
   wire \MEM[3][3] ;
   wire \MEM[3][2] ;
   wire \MEM[3][1] ;
   wire \MEM[3][0] ;
   wire \MEM[2][7] ;
   wire \MEM[2][6] ;
   wire \MEM[2][5] ;
   wire \MEM[2][4] ;
   wire \MEM[2][3] ;
   wire \MEM[2][2] ;
   wire \MEM[2][1] ;
   wire \MEM[2][0] ;
   wire \MEM[1][7] ;
   wire \MEM[1][6] ;
   wire \MEM[1][5] ;
   wire \MEM[1][4] ;
   wire \MEM[1][3] ;
   wire \MEM[1][2] ;
   wire \MEM[1][1] ;
   wire \MEM[1][0] ;
   wire \MEM[0][7] ;
   wire \MEM[0][6] ;
   wire \MEM[0][5] ;
   wire \MEM[0][4] ;
   wire \MEM[0][3] ;
   wire \MEM[0][2] ;
   wire \MEM[0][1] ;
   wire \MEM[0][0] ;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;

   assign N9 = raddr[0] ;
   assign N10 = raddr[1] ;
   assign N11 = raddr[2] ;
   assign test_so = \MEM[7][7]  ;

   // Module instantiations
   SDFFRQX2M \MEM_reg[5][7]  (
	.SI(\MEM[5][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[5][7] ),
	.D(n133),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][6]  (
	.SI(\MEM[5][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[5][6] ),
	.D(n132),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][5]  (
	.SI(\MEM[5][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[5][5] ),
	.D(n131),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][4]  (
	.SI(\MEM[5][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[5][4] ),
	.D(n130),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][3]  (
	.SI(\MEM[5][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[5][3] ),
	.D(n129),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][2]  (
	.SI(\MEM[5][1] ),
	.SE(n186),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[5][2] ),
	.D(n128),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][1]  (
	.SI(\MEM[5][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[5][1] ),
	.D(n127),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[5][0]  (
	.SI(\MEM[4][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[5][0] ),
	.D(n126),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][7]  (
	.SI(\MEM[1][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[1][7] ),
	.D(n101),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][6]  (
	.SI(\MEM[1][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[1][6] ),
	.D(n100),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][5]  (
	.SI(\MEM[1][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[1][5] ),
	.D(n99),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][4]  (
	.SI(\MEM[1][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[1][4] ),
	.D(n98),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][3]  (
	.SI(\MEM[1][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[1][3] ),
	.D(n97),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][2]  (
	.SI(\MEM[1][1] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[1][2] ),
	.D(n96),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][1]  (
	.SI(\MEM[1][0] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[1][1] ),
	.D(n95),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[1][0]  (
	.SI(\MEM[0][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[1][0] ),
	.D(n94),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][7]  (
	.SI(\MEM[7][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[7][7] ),
	.D(n149),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][6]  (
	.SI(\MEM[7][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[7][6] ),
	.D(n148),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][5]  (
	.SI(\MEM[7][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[7][5] ),
	.D(n147),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][4]  (
	.SI(\MEM[7][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[7][4] ),
	.D(n146),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][3]  (
	.SI(\MEM[7][2] ),
	.SE(n187),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[7][3] ),
	.D(n145),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][2]  (
	.SI(\MEM[7][1] ),
	.SE(n186),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[7][2] ),
	.D(n144),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][1]  (
	.SI(\MEM[7][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[7][1] ),
	.D(n143),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[7][0]  (
	.SI(\MEM[6][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[7][0] ),
	.D(n142),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][7]  (
	.SI(\MEM[3][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[3][7] ),
	.D(n117),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][6]  (
	.SI(\MEM[3][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[3][6] ),
	.D(n116),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][5]  (
	.SI(\MEM[3][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[3][5] ),
	.D(n115),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][4]  (
	.SI(\MEM[3][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[3][4] ),
	.D(n114),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][3]  (
	.SI(\MEM[3][2] ),
	.SE(n187),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[3][3] ),
	.D(n113),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][2]  (
	.SI(\MEM[3][1] ),
	.SE(n186),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[3][2] ),
	.D(n112),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][1]  (
	.SI(\MEM[3][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[3][1] ),
	.D(n111),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[3][0]  (
	.SI(\MEM[2][7] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[3][0] ),
	.D(n110),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][7]  (
	.SI(\MEM[6][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[6][7] ),
	.D(n141),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][6]  (
	.SI(\MEM[6][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[6][6] ),
	.D(n140),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][5]  (
	.SI(\MEM[6][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[6][5] ),
	.D(n139),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][4]  (
	.SI(\MEM[6][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[6][4] ),
	.D(n138),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][3]  (
	.SI(\MEM[6][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[6][3] ),
	.D(n137),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][2]  (
	.SI(\MEM[6][1] ),
	.SE(n186),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[6][2] ),
	.D(n136),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][1]  (
	.SI(\MEM[6][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[6][1] ),
	.D(n135),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[6][0]  (
	.SI(\MEM[5][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[6][0] ),
	.D(n134),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][7]  (
	.SI(\MEM[2][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[2][7] ),
	.D(n109),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][6]  (
	.SI(\MEM[2][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[2][6] ),
	.D(n108),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][5]  (
	.SI(\MEM[2][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[2][5] ),
	.D(n107),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][4]  (
	.SI(\MEM[2][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[2][4] ),
	.D(n106),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][3]  (
	.SI(\MEM[2][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[2][3] ),
	.D(n105),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][2]  (
	.SI(\MEM[2][1] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[2][2] ),
	.D(n104),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][1]  (
	.SI(\MEM[2][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[2][1] ),
	.D(n103),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[2][0]  (
	.SI(\MEM[1][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[2][0] ),
	.D(n102),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][7]  (
	.SI(\MEM[4][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[4][7] ),
	.D(n125),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][6]  (
	.SI(\MEM[4][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[4][6] ),
	.D(n124),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][5]  (
	.SI(\MEM[4][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[4][5] ),
	.D(n123),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][4]  (
	.SI(\MEM[4][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[4][4] ),
	.D(n122),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][3]  (
	.SI(\MEM[4][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[4][3] ),
	.D(n121),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][2]  (
	.SI(\MEM[4][1] ),
	.SE(n186),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[4][2] ),
	.D(n120),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][1]  (
	.SI(\MEM[4][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[4][1] ),
	.D(n119),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[4][0]  (
	.SI(\MEM[3][7] ),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[4][0] ),
	.D(n118),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][7]  (
	.SI(\MEM[0][6] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[0][7] ),
	.D(n93),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][6]  (
	.SI(\MEM[0][5] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[0][6] ),
	.D(n92),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][5]  (
	.SI(\MEM[0][4] ),
	.SE(n185),
	.RN(wrst_n),
	.Q(\MEM[0][5] ),
	.D(n91),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][4]  (
	.SI(\MEM[0][3] ),
	.SE(n184),
	.RN(wrst_n),
	.Q(\MEM[0][4] ),
	.D(n90),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][3]  (
	.SI(\MEM[0][2] ),
	.SE(n187),
	.RN(wrst_n),
	.Q(\MEM[0][3] ),
	.D(n89),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][2]  (
	.SI(\MEM[0][1] ),
	.SE(n186),
	.RN(wrst_n),
	.Q(\MEM[0][2] ),
	.D(n88),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][1]  (
	.SI(\MEM[0][0] ),
	.SE(n185),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[0][1] ),
	.D(n87),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \MEM_reg[0][0]  (
	.SI(test_si),
	.SE(n184),
	.RN(FE_OFN0_SYNC_REF_RST_M),
	.Q(\MEM[0][0] ),
	.D(n86),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U77 (
	.Y(n81),
	.C(n82),
	.B(n180),
	.A(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U78 (
	.Y(n75),
	.C(n76),
	.B(n180),
	.A(n179), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U79 (
	.Y(n80),
	.B(wfull),
	.AN(winc), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U80 (
	.Y(n79),
	.C(waddr[1]),
	.B(n76),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U81 (
	.Y(n76),
	.B(waddr[2]),
	.AN(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U82 (
	.Y(n86),
	.B1(n178),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n87),
	.B1(n177),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n88),
	.B1(n176),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n89),
	.B1(n175),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n90),
	.B1(n174),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n91),
	.B1(n173),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n92),
	.B1(n172),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n93),
	.B1(n171),
	.B0(n75),
	.A1N(n75),
	.A0N(\MEM[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n110),
	.B1(n79),
	.B0(n178),
	.A1N(n79),
	.A0N(\MEM[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n111),
	.B1(n79),
	.B0(n177),
	.A1N(n79),
	.A0N(\MEM[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n112),
	.B1(n79),
	.B0(n176),
	.A1N(n79),
	.A0N(\MEM[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n113),
	.B1(n79),
	.B0(n175),
	.A1N(n79),
	.A0N(\MEM[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n114),
	.B1(n79),
	.B0(n174),
	.A1N(n79),
	.A0N(\MEM[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n115),
	.B1(n79),
	.B0(n173),
	.A1N(n79),
	.A0N(\MEM[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n116),
	.B1(n79),
	.B0(n172),
	.A1N(n79),
	.A0N(\MEM[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n117),
	.B1(n79),
	.B0(n171),
	.A1N(n79),
	.A0N(\MEM[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n118),
	.B1(n81),
	.B0(n178),
	.A1N(n81),
	.A0N(\MEM[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n119),
	.B1(n81),
	.B0(n177),
	.A1N(n81),
	.A0N(\MEM[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n120),
	.B1(n81),
	.B0(n176),
	.A1N(n81),
	.A0N(\MEM[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n121),
	.B1(n81),
	.B0(n175),
	.A1N(n81),
	.A0N(\MEM[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n122),
	.B1(n81),
	.B0(n174),
	.A1N(n81),
	.A0N(\MEM[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n123),
	.B1(n81),
	.B0(n173),
	.A1N(n81),
	.A0N(\MEM[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n124),
	.B1(n81),
	.B0(n172),
	.A1N(n81),
	.A0N(\MEM[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n125),
	.B1(n81),
	.B0(n171),
	.A1N(n81),
	.A0N(\MEM[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n178),
	.A(wdata[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n177),
	.A(wdata[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n176),
	.A(wdata[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n175),
	.A(wdata[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U110 (
	.Y(n174),
	.A(wdata[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U111 (
	.Y(n173),
	.A(wdata[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U112 (
	.Y(n172),
	.A(wdata[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n171),
	.A(wdata[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U115 (
	.Y(n84),
	.C(n82),
	.B(n179),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U117 (
	.Y(n85),
	.C(n82),
	.B(waddr[0]),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n94),
	.B1(n77),
	.B0(n178),
	.A1N(n77),
	.A0N(\MEM[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n95),
	.B1(n77),
	.B0(n177),
	.A1N(n77),
	.A0N(\MEM[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n96),
	.B1(n77),
	.B0(n176),
	.A1N(n77),
	.A0N(\MEM[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n97),
	.B1(n77),
	.B0(n175),
	.A1N(n77),
	.A0N(\MEM[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n98),
	.B1(n77),
	.B0(n174),
	.A1N(n77),
	.A0N(\MEM[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n99),
	.B1(n77),
	.B0(n173),
	.A1N(n77),
	.A0N(\MEM[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n100),
	.B1(n77),
	.B0(n172),
	.A1N(n77),
	.A0N(\MEM[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n101),
	.B1(n77),
	.B0(n171),
	.A1N(n77),
	.A0N(\MEM[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n102),
	.B1(n78),
	.B0(n178),
	.A1N(n78),
	.A0N(\MEM[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U127 (
	.Y(n103),
	.B1(n78),
	.B0(n177),
	.A1N(n78),
	.A0N(\MEM[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U128 (
	.Y(n104),
	.B1(n78),
	.B0(n176),
	.A1N(n78),
	.A0N(\MEM[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U129 (
	.Y(n105),
	.B1(n78),
	.B0(n175),
	.A1N(n78),
	.A0N(\MEM[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U130 (
	.Y(n106),
	.B1(n78),
	.B0(n174),
	.A1N(n78),
	.A0N(\MEM[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U131 (
	.Y(n107),
	.B1(n78),
	.B0(n173),
	.A1N(n78),
	.A0N(\MEM[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U132 (
	.Y(n108),
	.B1(n78),
	.B0(n172),
	.A1N(n78),
	.A0N(\MEM[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U133 (
	.Y(n109),
	.B1(n78),
	.B0(n171),
	.A1N(n78),
	.A0N(\MEM[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U134 (
	.Y(n126),
	.B1(n83),
	.B0(n178),
	.A1N(n83),
	.A0N(\MEM[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U135 (
	.Y(n127),
	.B1(n83),
	.B0(n177),
	.A1N(n83),
	.A0N(\MEM[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n128),
	.B1(n83),
	.B0(n176),
	.A1N(n83),
	.A0N(\MEM[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n129),
	.B1(n83),
	.B0(n175),
	.A1N(n83),
	.A0N(\MEM[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n130),
	.B1(n83),
	.B0(n174),
	.A1N(n83),
	.A0N(\MEM[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n131),
	.B1(n83),
	.B0(n173),
	.A1N(n83),
	.A0N(\MEM[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n132),
	.B1(n83),
	.B0(n172),
	.A1N(n83),
	.A0N(\MEM[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n133),
	.B1(n83),
	.B0(n171),
	.A1N(n83),
	.A0N(\MEM[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n134),
	.B1(n84),
	.B0(n178),
	.A1N(n84),
	.A0N(\MEM[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n135),
	.B1(n84),
	.B0(n177),
	.A1N(n84),
	.A0N(\MEM[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n136),
	.B1(n84),
	.B0(n176),
	.A1N(n84),
	.A0N(\MEM[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n137),
	.B1(n84),
	.B0(n175),
	.A1N(n84),
	.A0N(\MEM[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n138),
	.B1(n84),
	.B0(n174),
	.A1N(n84),
	.A0N(\MEM[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n139),
	.B1(n84),
	.B0(n173),
	.A1N(n84),
	.A0N(\MEM[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n140),
	.B1(n84),
	.B0(n172),
	.A1N(n84),
	.A0N(\MEM[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U149 (
	.Y(n141),
	.B1(n84),
	.B0(n171),
	.A1N(n84),
	.A0N(\MEM[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U150 (
	.Y(n142),
	.B1(n85),
	.B0(n178),
	.A1N(n85),
	.A0N(\MEM[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U151 (
	.Y(n143),
	.B1(n85),
	.B0(n177),
	.A1N(n85),
	.A0N(\MEM[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U152 (
	.Y(n144),
	.B1(n85),
	.B0(n176),
	.A1N(n85),
	.A0N(\MEM[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U153 (
	.Y(n145),
	.B1(n85),
	.B0(n175),
	.A1N(n85),
	.A0N(\MEM[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U154 (
	.Y(n146),
	.B1(n85),
	.B0(n174),
	.A1N(n85),
	.A0N(\MEM[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U155 (
	.Y(n147),
	.B1(n85),
	.B0(n173),
	.A1N(n85),
	.A0N(\MEM[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U156 (
	.Y(n148),
	.B1(n85),
	.B0(n172),
	.A1N(n85),
	.A0N(\MEM[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U157 (
	.Y(n149),
	.B1(n85),
	.B0(n171),
	.A1N(n85),
	.A0N(\MEM[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U158 (
	.Y(n83),
	.C(n82),
	.B(n180),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U159 (
	.Y(n82),
	.B(n80),
	.A(waddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U160 (
	.Y(n78),
	.C(waddr[1]),
	.B(n179),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U161 (
	.Y(n77),
	.C(waddr[0]),
	.B(n180),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U162 (
	.Y(n180),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U163 (
	.Y(n179),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U164 (
	.Y(rdata[6]),
	.S0(N11),
	.B(n152),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U165 (
	.Y(n153),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][6] ),
	.C(\MEM[2][6] ),
	.B(\MEM[1][6] ),
	.A(\MEM[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U166 (
	.Y(n152),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][6] ),
	.C(\MEM[6][6] ),
	.B(\MEM[5][6] ),
	.A(\MEM[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U167 (
	.Y(rdata[7]),
	.S0(N11),
	.B(n154),
	.A(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U168 (
	.Y(n155),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][7] ),
	.C(\MEM[2][7] ),
	.B(\MEM[1][7] ),
	.A(\MEM[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U169 (
	.Y(n154),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][7] ),
	.C(\MEM[6][7] ),
	.B(\MEM[5][7] ),
	.A(\MEM[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U170 (
	.Y(rdata[3]),
	.S0(N11),
	.B(n71),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U171 (
	.Y(n72),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][3] ),
	.C(\MEM[2][3] ),
	.B(\MEM[1][3] ),
	.A(\MEM[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U172 (
	.Y(n71),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][3] ),
	.C(\MEM[6][3] ),
	.B(\MEM[5][3] ),
	.A(\MEM[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U173 (
	.Y(rdata[4]),
	.S0(N11),
	.B(n73),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U174 (
	.Y(n74),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][4] ),
	.C(\MEM[2][4] ),
	.B(\MEM[1][4] ),
	.A(\MEM[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U175 (
	.Y(n73),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][4] ),
	.C(\MEM[6][4] ),
	.B(\MEM[5][4] ),
	.A(\MEM[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U176 (
	.Y(rdata[0]),
	.S0(N11),
	.B(n65),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U177 (
	.Y(n66),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][0] ),
	.C(\MEM[2][0] ),
	.B(\MEM[1][0] ),
	.A(\MEM[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U178 (
	.Y(n65),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][0] ),
	.C(\MEM[6][0] ),
	.B(\MEM[5][0] ),
	.A(\MEM[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U179 (
	.Y(rdata[5]),
	.S0(N11),
	.B(n150),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U180 (
	.Y(n151),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][5] ),
	.C(\MEM[2][5] ),
	.B(\MEM[1][5] ),
	.A(\MEM[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U181 (
	.Y(n150),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][5] ),
	.C(\MEM[6][5] ),
	.B(\MEM[5][5] ),
	.A(\MEM[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U182 (
	.Y(rdata[1]),
	.S0(N11),
	.B(n67),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U183 (
	.Y(n68),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][1] ),
	.C(\MEM[2][1] ),
	.B(\MEM[1][1] ),
	.A(\MEM[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U184 (
	.Y(n67),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][1] ),
	.C(\MEM[6][1] ),
	.B(\MEM[5][1] ),
	.A(\MEM[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U185 (
	.Y(rdata[2]),
	.S0(N11),
	.B(n69),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U186 (
	.Y(n70),
	.S1(N10),
	.S0(n157),
	.D(\MEM[3][2] ),
	.C(\MEM[2][2] ),
	.B(\MEM[1][2] ),
	.A(\MEM[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U187 (
	.Y(n69),
	.S1(N10),
	.S0(n156),
	.D(\MEM[7][2] ),
	.C(\MEM[6][2] ),
	.B(\MEM[5][2] ),
	.A(\MEM[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U188 (
	.Y(n156),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U189 (
	.Y(n157),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U190 (
	.Y(n183),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U191 (
	.Y(n184),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U192 (
	.Y(n185),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U193 (
	.Y(n186),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U194 (
	.Y(n187),
	.A(n183), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module r_empty_P_SIZE4_test_1 (
	rinc, 
	rclk, 
	rrst_n, 
	rq2_wptr, 
	rempty, 
	raddr, 
	g_rptr, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input rinc;
   input rclk;
   input rrst_n;
   input [3:0] rq2_wptr;
   output rempty;
   output [2:0] raddr;
   output [3:0] g_rptr;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \bn_rptr[3] ;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n1;
   wire n2;
   wire n11;
   wire n12;

   // Module instantiations
   SDFFRQX2M \g_rptr_reg[0]  (
	.SI(n12),
	.SE(test_se),
	.RN(rrst_n),
	.Q(g_rptr[0]),
	.D(n41),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_rptr_reg[3]  (
	.SI(g_rptr[2]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(g_rptr[3]),
	.D(n34),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_rptr_reg[2]  (
	.SI(g_rptr[1]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(g_rptr[2]),
	.D(n35),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_rptr_reg[1]  (
	.SI(g_rptr[0]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(g_rptr[1]),
	.D(n36),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_rptr_reg[3]  (
	.SI(n11),
	.SE(test_se),
	.RN(rrst_n),
	.Q(\bn_rptr[3] ),
	.D(n37),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_rptr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddr[0]),
	.D(n40),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_rptr_reg[2]  (
	.SI(n2),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddr[2]),
	.D(n38),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \bn_rptr_reg[1]  (
	.SI(raddr[0]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddr[1]),
	.D(n39),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U11 (
	.Y(n16),
	.C(n17),
	.B(n2),
	.AN(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(n21),
	.B1(n19),
	.B0(n2),
	.A1N(n24),
	.A0N(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U13 (
	.Y(n39),
	.B(n27),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n32),
	.B(rq2_wptr[2]),
	.A(g_rptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U16 (
	.Y(n17),
	.C0(n19),
	.B0(n22),
	.A1(n12),
	.A0(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U17 (
	.Y(n38),
	.B(n26),
	.A(raddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U18 (
	.Y(n27),
	.B(n28),
	.AN(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n40),
	.B(n28),
	.A(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U20 (
	.Y(rempty),
	.D(n32),
	.C(n31),
	.B(n30),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U21 (
	.Y(n29),
	.B(rq2_wptr[1]),
	.A(g_rptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U22 (
	.Y(n30),
	.B(rq2_wptr[0]),
	.A(g_rptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U23 (
	.Y(n31),
	.B(rq2_wptr[3]),
	.A(g_rptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U24 (
	.Y(n37),
	.C0(n19),
	.B0(n25),
	.A1(n12),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U25 (
	.Y(n25),
	.C(n1),
	.B(n12),
	.A(raddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n1),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U27 (
	.Y(n35),
	.C0(n20),
	.B0(n19),
	.A1(n18),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U28 (
	.Y(n20),
	.B0(n21),
	.A1(g_rptr[2]),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U29 (
	.Y(n36),
	.C0(n23),
	.B0(n22),
	.A1(n18),
	.A0(raddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U30 (
	.Y(n23),
	.B0(n21),
	.A1(g_rptr[1]),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(n24),
	.B(raddr[1]),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n18),
	.B(n12),
	.A(raddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U33 (
	.Y(n26),
	.B(raddr[1]),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U34 (
	.Y(n19),
	.B(n11),
	.A(\bn_rptr[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U35 (
	.Y(n2),
	.A(raddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n11),
	.A(raddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n12),
	.A(\bn_rptr[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(n28),
	.B(rempty),
	.A(rinc), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U39 (
	.Y(n22),
	.B(\bn_rptr[3] ),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U40 (
	.Y(n41),
	.B0(n33),
	.A1N(n16),
	.A0N(g_rptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U41 (
	.Y(n33),
	.B(raddr[1]),
	.A(raddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U42 (
	.Y(n34),
	.B0(n17),
	.A1(n16),
	.A0(g_rptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module w_full_POI_SIZE4_test_1 (
	winc, 
	wclk, 
	wrst_n, 
	wq2_rptr, 
	wfull, 
	waddr, 
	g_wptr, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input winc;
   input wclk;
   input wrst_n;
   input [3:0] wq2_rptr;
   output wfull;
   output [2:0] waddr;
   output [3:0] g_wptr;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \bn_wptr[3] ;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n1;
   wire n2;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;

   // Module instantiations
   SDFFRQX2M \g_wptr_reg[3]  (
	.SI(g_wptr[2]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(g_wptr[3]),
	.D(n39),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_wptr_reg[0]  (
	.SI(n15),
	.SE(test_se),
	.RN(wrst_n),
	.Q(g_wptr[0]),
	.D(n1),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_wptr_reg[1]  (
	.SI(g_wptr[0]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(g_wptr[1]),
	.D(n12),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \g_wptr_reg[2]  (
	.SI(g_wptr[1]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(g_wptr[2]),
	.D(n40),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_wptr_reg[3]  (
	.SI(waddr[2]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(\bn_wptr[3] ),
	.D(n41),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_wptr_reg[2]  (
	.SI(n13),
	.SE(test_se),
	.RN(wrst_n),
	.Q(waddr[2]),
	.D(n42),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_wptr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(wrst_n),
	.Q(waddr[0]),
	.D(n44),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bn_wptr_reg[1]  (
	.SI(n11),
	.SE(test_se),
	.RN(wrst_n),
	.Q(waddr[1]),
	.D(n43),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U11 (
	.Y(n20),
	.C0(n22),
	.B0(n27),
	.A1N(n38),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U12 (
	.Y(n19),
	.C(n20),
	.B(n24),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U13 (
	.Y(n43),
	.B(n31),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n32),
	.B(n18),
	.A(winc), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(wfull),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(n21),
	.B(n15),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U17 (
	.Y(n35),
	.B(n15),
	.A(g_wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(n28),
	.B(waddr[1]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n44),
	.B(n32),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U20 (
	.Y(n42),
	.B(n30),
	.A(waddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n13),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(n31),
	.B(n11),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n11),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U24 (
	.Y(n18),
	.D(n36),
	.C(n35),
	.B(n34),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U25 (
	.Y(n36),
	.B(g_wptr[2]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U26 (
	.Y(n33),
	.B(waddr[0]),
	.A(g_wptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U27 (
	.Y(n34),
	.B(waddr[1]),
	.A(g_wptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U28 (
	.Y(n41),
	.C0(n22),
	.B0(n29),
	.A1(n15),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U29 (
	.Y(n29),
	.C(n2),
	.B(n15),
	.A(waddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n2),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n30),
	.B(waddr[1]),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n15),
	.A(\bn_wptr[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(n38),
	.B(waddr[0]),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n14),
	.A(waddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U35 (
	.Y(n27),
	.B(\bn_wptr[3] ),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n1),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U37 (
	.Y(n37),
	.C0(n38),
	.B1(n19),
	.B0(g_wptr[0]),
	.A1(waddr[0]),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n12),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U39 (
	.Y(n25),
	.C0(n26),
	.B1(n19),
	.B0(g_wptr[1]),
	.A1(n24),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U40 (
	.Y(n26),
	.C0(n27),
	.B0(n21),
	.A1(n13),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U41 (
	.Y(n40),
	.C(n23),
	.B(n22),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U42 (
	.Y(n23),
	.B1(g_wptr[2]),
	.B0(n19),
	.A1(waddr[2]),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U43 (
	.Y(n39),
	.B0(n20),
	.A1(n19),
	.A0(g_wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U44 (
	.Y(n24),
	.B(\bn_wptr[3] ),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U45 (
	.Y(n22),
	.B(n14),
	.A(\bn_wptr[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_CTRL_test_1 (
	RX_P_DATA, 
	RX_D_VLD, 
	FIFO_FULL, 
	ALU_OUT, 
	OUT_Valid, 
	Rd_D_Vld, 
	Rd_D, 
	CLK, 
	RST, 
	WR_DATA, 
	WR_INC, 
	ALU_EN, 
	ALU_FUN, 
	Wr_D, 
	Addr, 
	RdEn, 
	CLK_EN, 
	CLK_DIV_EN, 
	WrEn, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] RX_P_DATA;
   input RX_D_VLD;
   input FIFO_FULL;
   input [15:0] ALU_OUT;
   input OUT_Valid;
   input Rd_D_Vld;
   input [7:0] Rd_D;
   input CLK;
   input RST;
   output [7:0] WR_DATA;
   output WR_INC;
   output ALU_EN;
   output [3:0] ALU_FUN;
   output [7:0] Wr_D;
   output [3:0] Addr;
   output RdEn;
   output CLK_EN;
   output CLK_DIV_EN;
   output WrEn;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n64;
   wire n65;
   wire n66;
   wire [3:0] current_state;
   wire [3:0] next_state;

   assign test_so = n16 ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(n18),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[3]),
	.D(next_state[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n11),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(Addr[1]),
	.B(n64),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(ALU_FUN[2]),
	.B(n12),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n12),
	.A(ALU_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(WrEn),
	.B(n39),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(ALU_EN),
	.B(n42),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U16 (
	.Y(n51),
	.B0(n27),
	.A1(n66),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(ALU_FUN[3]),
	.B(n12),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(ALU_FUN[0]),
	.B(n12),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(Addr[0]),
	.B(n40),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U20 (
	.Y(ALU_FUN[1]),
	.B(n12),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U21 (
	.Y(n24),
	.B(n30),
	.AN(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(Addr[2]),
	.B(n40),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(Wr_D[5]),
	.B(n19),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(Wr_D[1]),
	.B(n64),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(Wr_D[2]),
	.B(n22),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(Wr_D[3]),
	.B(n21),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U27 (
	.Y(Wr_D[4]),
	.B(n20),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U28 (
	.Y(Wr_D[0]),
	.B(n65),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U29 (
	.Y(n39),
	.B(n16),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n9),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(Addr[3]),
	.B(n40),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n27),
	.B(n52),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(RdEn),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n15),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U35 (
	.Y(n14),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n10),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U37 (
	.Y(n52),
	.B(current_state[3]),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n42),
	.C(current_state[2]),
	.B(n52),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n17),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U40 (
	.Y(n30),
	.C(n18),
	.B(current_state[0]),
	.AN(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U41 (
	.Y(n53),
	.C(n18),
	.B(current_state[3]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U42 (
	.Y(n40),
	.C(current_state[0]),
	.B(n18),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U43 (
	.Y(n33),
	.B(current_state[0]),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n65),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n64),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n22),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n18),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n66),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n21),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U50 (
	.Y(WR_INC),
	.C0(n55),
	.B0(n54),
	.A1N(OUT_Valid),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U51 (
	.Y(n32),
	.C(n11),
	.B(current_state[2]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U52 (
	.Y(n34),
	.C0(n23),
	.B0(n41),
	.A1(n40),
	.A0(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U53 (
	.Y(n41),
	.C(n46),
	.B(RX_P_DATA[0]),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U54 (
	.Y(n49),
	.B(current_state[0]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U55 (
	.Y(n54),
	.D(n53),
	.C(Rd_D_Vld),
	.B(n11),
	.AN(FIFO_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U56 (
	.Y(Wr_D[6]),
	.B(n51),
	.AN(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U57 (
	.Y(Wr_D[7]),
	.B(n51),
	.AN(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U58 (
	.Y(next_state[1]),
	.C0(n28),
	.B0(n13),
	.A1(n27),
	.A0(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U59 (
	.Y(n28),
	.C0(n30),
	.B0(n10),
	.A1(n29),
	.A0(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U60 (
	.Y(n13),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U61 (
	.Y(n29),
	.B(n33),
	.AN(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U62 (
	.Y(n55),
	.D(current_state[3]),
	.C(current_state[1]),
	.B(n49),
	.A(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U63 (
	.Y(n45),
	.D(n50),
	.C(RX_P_DATA[7]),
	.B(n49),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U64 (
	.Y(n50),
	.C(current_state[1]),
	.B(current_state[3]),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U65 (
	.Y(n63),
	.B1(n15),
	.B0(ALU_OUT[8]),
	.A1(n9),
	.A0(Rd_D[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U66 (
	.Y(n31),
	.B(current_state[3]),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U67 (
	.Y(WR_DATA[1]),
	.B0(n62),
	.A1N(n14),
	.A0N(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U68 (
	.Y(n62),
	.B1(n15),
	.B0(ALU_OUT[9]),
	.A1(n9),
	.A0(Rd_D[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U69 (
	.Y(WR_DATA[2]),
	.B0(n61),
	.A1N(n14),
	.A0N(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U70 (
	.Y(n61),
	.B1(n15),
	.B0(ALU_OUT[10]),
	.A1(n9),
	.A0(Rd_D[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U71 (
	.Y(WR_DATA[3]),
	.B0(n60),
	.A1N(n14),
	.A0N(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U72 (
	.Y(n60),
	.B1(n15),
	.B0(ALU_OUT[11]),
	.A1(n9),
	.A0(Rd_D[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U73 (
	.Y(WR_DATA[4]),
	.B0(n59),
	.A1N(n14),
	.A0N(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U74 (
	.Y(n59),
	.B1(n15),
	.B0(ALU_OUT[12]),
	.A1(n9),
	.A0(Rd_D[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U75 (
	.Y(WR_DATA[5]),
	.B0(n58),
	.A1N(n14),
	.A0N(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U76 (
	.Y(n58),
	.B1(n15),
	.B0(ALU_OUT[13]),
	.A1(n9),
	.A0(Rd_D[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U77 (
	.Y(WR_DATA[6]),
	.B0(n57),
	.A1N(n14),
	.A0N(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U78 (
	.Y(n57),
	.B1(n15),
	.B0(ALU_OUT[14]),
	.A1(n9),
	.A0(Rd_D[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U79 (
	.Y(WR_DATA[7]),
	.B0(n56),
	.A1N(n14),
	.A0N(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U80 (
	.Y(n56),
	.B1(n15),
	.B0(ALU_OUT[15]),
	.A1(n9),
	.A0(Rd_D[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U81 (
	.Y(n46),
	.D(n45),
	.C(n47),
	.B(RX_P_DATA[1]),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U82 (
	.Y(n47),
	.B(RX_P_DATA[2]),
	.A(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA22X2M U83 (
	.Y(n23),
	.B1(n44),
	.B0(n43),
	.A1(n42),
	.A0(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U84 (
	.Y(n44),
	.C(RX_P_DATA[4]),
	.B(RX_P_DATA[6]),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U85 (
	.Y(n43),
	.D(n19),
	.C(n64),
	.B(n45),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U86 (
	.Y(next_state[0]),
	.D(n37),
	.C(n36),
	.B(n26),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U87 (
	.Y(n36),
	.C(n46),
	.B(n20),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U88 (
	.Y(n37),
	.C0(n38),
	.B0(n34),
	.A1(RX_D_VLD),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U89 (
	.Y(n38),
	.B0(RX_D_VLD),
	.A1(n39),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U90 (
	.Y(n16),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U91 (
	.Y(n11),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U92 (
	.Y(next_state[3]),
	.B0(n12),
	.A2(current_state[1]),
	.A1(current_state[2]),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U93 (
	.Y(n35),
	.D(n17),
	.C(current_state[3]),
	.B(n49),
	.A(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U94 (
	.Y(n26),
	.D(n48),
	.C(RX_P_DATA[6]),
	.B(n45),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U95 (
	.Y(n48),
	.D(RX_P_DATA[0]),
	.C(RX_P_DATA[1]),
	.B(RX_P_DATA[4]),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U96 (
	.Y(n20),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n19),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U98 (
	.Y(next_state[2]),
	.C(n25),
	.B(n24),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U99 (
	.Y(n25),
	.B0N(n26),
	.A1(RX_D_VLD),
	.A0(RdEn), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U100 (
	.Y(WR_DATA[0]),
	.B0(n63),
	.A1N(n14),
	.A0N(ALU_OUT[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(CLK_DIV_EN),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(CLK_EN),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Pulse_Gen_test_1 (
	CLK, 
	RST, 
	en_sig, 
	Pulse_en, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input en_sig;
   output Pulse_en;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire sync_flop;
   wire meta_flop;

   assign test_so = sync_flop ;

   // Module instantiations
   SDFFRQX2M meta_flop_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(meta_flop),
	.D(en_sig),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M sync_flop_reg (
	.SI(meta_flop),
	.SE(test_se),
	.RN(RST),
	.Q(sync_flop),
	.D(meta_flop),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U6 (
	.Y(Pulse_en),
	.B(sync_flop),
	.AN(meta_flop), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYSTEM (
	REF_CLK, 
	RST, 
	UART_CLK, 
	UART_RX_IN, 
	scan_clk, 
	scan_reset, 
	test_mode, 
	SE, 
	SI, 
	SO, 
	UART_TX_OUT, 
	VDD, 
	VSS);
   input REF_CLK;
   input RST;
   input UART_CLK;
   input UART_RX_IN;
   input scan_clk;
   input scan_reset;
   input test_mode;
   input SE;
   input [3:0] SI;
   output [3:0] SO;
   output UART_TX_OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N1;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire REF_CLK_M__L2_N1;
   wire REF_CLK_M__L2_N0;
   wire REF_CLK_M__L1_N0;
   wire UART_CLK_M__L7_N1;
   wire UART_CLK_M__L7_N0;
   wire UART_CLK_M__L6_N2;
   wire UART_CLK_M__L6_N1;
   wire UART_CLK_M__L6_N0;
   wire UART_CLK_M__L5_N1;
   wire UART_CLK_M__L5_N0;
   wire UART_CLK_M__L4_N1;
   wire UART_CLK_M__L4_N0;
   wire UART_CLK_M__L3_N1;
   wire UART_CLK_M__L3_N0;
   wire UART_CLK_M__L2_N3;
   wire UART_CLK_M__L2_N2;
   wire UART_CLK_M__L2_N1;
   wire UART_CLK_M__L2_N0;
   wire UART_CLK_M__L1_N1;
   wire UART_CLK_M__L1_N0;
   wire UART_TX_CLK_M__L1_N0;
   wire UART_RX_CLK_M__L1_N0;
   wire FE_OFN4_SE;
   wire FE_OFN3_SYNC_UART_RST_M;
   wire FE_OFN0_SYNC_REF_RST_M;
   wire REF_CLK_M;
   wire UART_CLK_M;
   wire RST_M;
   wire SYNC_REF_RST;
   wire SYNC_REF_RST_M;
   wire SYNC_UART_RST;
   wire SYNC_UART_RST_M;
   wire UART_RX_Vld_OUT;
   wire UART_RX_Vld_SYNC;
   wire UART_TX_CLK;
   wire UART_TX_CLK_M;
   wire UART_RX_CLK;
   wire UART_RX_CLK_M;
   wire _1_net_;
   wire ALU_CLK;
   wire RF_WrEn;
   wire RF_RdEn;
   wire RF_RdData_VLD;
   wire ALU_EN;
   wire ALU_OUT_VLD;
   wire UART_TX_Busy;
   wire F_EMPTY;
   wire WR_INC;
   wire RD_INC;
   wire FIFO_FULL;
   wire n2;
   wire n9;
   wire n10;
   wire n11;
   wire n15;
   wire n16;
   wire n17;
   wire n20;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire [7:0] UART_RX_OUT;
   wire [7:0] UART_RX_SYNC;
   wire [7:0] DIV_RATIO;
   wire [3:0] Addr;
   wire [7:0] Wr_D;
   wire [7:0] RF_RdData;
   wire [7:0] Op_A;
   wire [7:0] Op_B;
   wire [7:0] UART_Config;
   wire [3:0] ALU_FUN;
   wire [15:0] ALU_OUT;
   wire [7:0] RD_DATA;
   wire [7:0] WR_DATA;

   assign SO[2] = DIV_RATIO[2] ;
   assign _1_net_ = test_mode ;
endmodule

